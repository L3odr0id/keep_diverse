// Seed: 10701314730660828924,3128299129089410139

module zmouqukn
  (output byte hytib, input bit tjfijzhto [2:1][1:0], input logic on);
  
  
  not aeivfhvd(bqrt, jsf);
  
  nand tx(tg, on, on);
  
  or rx(hytib, hytib, tg);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic hytib -> byte hytib
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte hytib -> logic hytib
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jsf = 'b100zz;
  assign bqrt = 'b000;
  assign tg = 'b111;
endmodule: zmouqukn

module zcqb
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: zcqb

module pwurzywy
  (output logic [4:1][3:1] zaxcfri [4:2], input reg rjzcfsho, input triand logic [2:2][4:0] zhaane [3:3], input uwire logic xwbyuonkvi [2:1][2:4][2:3]);
  
  
  and yuwsigkms(bwcfnuxysf, bwcfnuxysf, bwcfnuxysf);
  
  not bynobzuy(bwcfnuxysf, bwcfnuxysf);
  
  
  // Single-driven assigns
  assign zaxcfri = '{'{'{'b0011x,'b1x1x1,'b0},'{'b0x,'b1,'bz},'{'b101zz,'bxz1,'b00x},'{'b00xz,'b00z01,'b01z}},'{'{'bx,'b1x,'b1},'{'bx1xxz,'b1,'bx0x},'{'bx1,'bx,'b00},'{'bxzxzz,'bz1xzz,'b11z}},'{'{'b0001,'b11,'b1},'{'b0,'b00x,'bzz},'{'b01,'b11,'b1zz0},'{'b1z00,'bz01z,'b0}}};
  
  // Multi-driven assigns
  assign zhaane = '{'{'{'b1x1,'b0,'bz1100,'bx1zz,'bzzx1z}}};
  assign bwcfnuxysf = 'b1z10;
endmodule: pwurzywy



// Seed after: 9741254061059762472,3128299129089410139
