// Seed: 2167559344450510339,3128299129089410139

module ybaupixgdc
  ( output wor logic [3:1][2:4] ytwms [0:0]
  , input tri0 logic yaphzgzxp [3:3]
  , input bit [2:3][3:3]  onqspnjr
  , input logic xlmgqjxv
  );
  
  
  not clgg(vapzajwwgt, onqspnjr);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][3:3]  onqspnjr -> logic onqspnjr
  
  or gcge(wqtvwavk, onqspnjr, wqtvwavk);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][3:3]  onqspnjr -> logic onqspnjr
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ybaupixgdc

module abwza
  (output reg [2:0][0:1]  cfsbpx, output reg lsf);
  
  wor logic [3:1][2:4] oeg [0:0];
  tri0 logic mzrljh [3:3];
  
  nand ubq(egekvrzt, hhtazbhdqq, ugw);
  
  ybaupixgdc uff(.ytwms(oeg), .yaphzgzxp(mzrljh), .onqspnjr(cfsbpx), .xlmgqjxv(cfsbpx));
  // warning: implicit conversion of port connection truncates from 6 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   reg [2:0][0:1]  cfsbpx -> bit [2:3][3:3]  onqspnjr
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   reg [2:0][0:1]  cfsbpx -> logic xlmgqjxv
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign egekvrzt = hhtazbhdqq;
  assign mzrljh = mzrljh;
endmodule: abwza

module g
  ( input wor logic [1:3][1:4] kydvey [2:4][2:1]
  , input trireg logic [1:3][4:4][3:0][2:4] zlllir [3:0][4:2]
  , input reg [2:3][0:2][0:3]  dc
  , input logic [0:4][0:4][0:3]  cgas
  );
  
  wor logic [3:1][2:4] ycwdqoabbe [0:0];
  wor logic [3:1][2:4] kwrigjfcxn [0:0];
  wor logic [3:1][2:4] flrzg [0:0];
  tri0 logic gqnhlcsa [3:3];
  tri0 logic nuxdgiypa [3:3];
  
  ybaupixgdc jgubwz(.ytwms(flrzg), .yaphzgzxp(nuxdgiypa), .onqspnjr(dc), .xlmgqjxv(dc));
  // warning: implicit conversion of port connection truncates from 24 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   reg [2:3][0:2][0:3]  dc -> bit [2:3][3:3]  onqspnjr
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   reg [2:3][0:2][0:3]  dc -> logic xlmgqjxv
  
  ybaupixgdc gbedgnsdat(.ytwms(kwrigjfcxn), .yaphzgzxp(nuxdgiypa), .onqspnjr(dc), .xlmgqjxv(s));
  // warning: implicit conversion of port connection truncates from 24 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   reg [2:3][0:2][0:3]  dc -> bit [2:3][3:3]  onqspnjr
  
  ybaupixgdc ganhf(.ytwms(ycwdqoabbe), .yaphzgzxp(gqnhlcsa), .onqspnjr(bk), .xlmgqjxv(s));
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic bk -> bit [2:3][3:3]  onqspnjr
  
  not qv(s, dc);
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   reg [2:3][0:2][0:3]  dc -> logic dc
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign gqnhlcsa = '{'b1x};
  assign nuxdgiypa = '{'bz};
  assign ycwdqoabbe = '{'{'{'b10xx,'b010,'bz},'{'b10,'bx100,'b0},'{'bx,'b11z0,'b011}}};
endmodule: g



// Seed after: 11767764356932420300,3128299129089410139
