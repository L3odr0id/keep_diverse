// Seed: 5290427713959618967,3128299129089410139

module fsxnq
  (output supply0 logic [0:1][2:4][3:2] piyauwq [0:1][1:3][3:0], input supply1 logic [4:4][0:3][2:4]  vwz);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign piyauwq = piyauwq;
endmodule: fsxnq

module jngnrxfen
  ();
  
  supply0 logic [0:1][2:4][3:2] jyefxedd [0:1][1:3][3:0];
  
  xor pu(t, t, hedc);
  
  and vmdupaf(t, hpcezcituq, ytsyiz);
  
  fsxnq fijvalhedk(.piyauwq(jyefxedd), .vwz(ouqoheom));
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic ouqoheom -> supply1 logic [4:4][0:3][2:4]  vwz
  
  and oytoxziav(c, wbcla, t);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign c = 'bx1x01;
  assign ytsyiz = t;
  assign hpcezcituq = hpcezcituq;
  assign hedc = 'b10z;
  assign t = t;
endmodule: jngnrxfen

module ag
  ( output shortreal totkrxnib [4:3]
  , output wand logic [3:0][3:1][3:3][1:3] cqvfp [4:4][3:3][3:1]
  , output byte qacaep [0:2]
  , output bit [0:0] v [4:2]
  );
  
  
  not abm(da, h);
  
  not dlkhctaycu(s, joy);
  
  or ddvtoijn(qzg, da, joy);
  
  
  // Single-driven assigns
  assign totkrxnib = totkrxnib;
  assign v = v;
  assign qacaep = '{'b0111,'b0111,'b00100};
  
  // Multi-driven assigns
  assign joy = 'bz01x0;
  assign da = 'bx0x;
  assign h = 'b0x0;
  assign cqvfp = cqvfp;
endmodule: ag

module htpzowxjx
  ( output logic [0:0][0:4][1:0][3:2]  ycf
  , input trior logic [3:4][3:3] orcan [2:0][1:0]
  , input supply1 logic [0:3][0:1][4:2][1:3] xjppsljm [1:2][3:4][0:2]
  , input triand logic [4:4][1:3][3:3]  aj
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: htpzowxjx



// Seed after: 16301470472216710936,3128299129089410139
