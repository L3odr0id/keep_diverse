// Seed: 8128931952326600637,3128299129089410139

module dhrf
  (output supply0 logic [2:1][1:4][4:1] nvgdrt [1:1][2:2], output bit [0:4][1:2][3:4]  mjoldlywo);
  
  
  
  // Single-driven assigns
  assign mjoldlywo = mjoldlywo;
  
  // Multi-driven assigns
  assign nvgdrt = nvgdrt;
endmodule: dhrf



// Seed after: 6823947585183604141,3128299129089410139
