// Seed: 16013029700436987217,3128299129089410139

module qgx
  ( output supply0 logic [0:4][2:3][1:1][2:4] dr [4:0][2:1][0:1]
  , input tri0 logic sz
  , input trior logic [4:1][1:3][2:4][3:4] vbptxvsm [4:3][4:0][2:0][2:0]
  , input tri0 logic [2:3][1:0] zvf [0:0][2:2][1:2]
  );
  
  
  not bdznex(ii, sz);
  
  xor xzyjmgu(iien, vmvuhyuhm, oakyqt);
  
  nand qxpuant(iien, sz, lyu);
  
  not ctp(lyu, mocr);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dr = dr;
  assign vmvuhyuhm = sz;
  assign oakyqt = 'b0;
  assign sz = 'bz1x;
  assign mocr = iien;
endmodule: qgx



// Seed after: 13278935458753096407,3128299129089410139
