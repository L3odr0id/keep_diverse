// Seed: 16397190719548895153,3128299129089410139

module tyiorvlgtp
  ( output logic [4:4][4:1]  dchlyvx
  , output bit [2:2][3:3] joojcolzhe [2:2]
  , output longint rztc
  , output wire logic [3:4][3:4][1:1] xdzgbddrf [3:0][3:2]
  , input wor logic xiphfxou [2:2][1:0][1:0][3:2]
  , input reg [0:0][1:3] dbgyjvigtf [4:1]
  , input bit [2:4]  i
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: tyiorvlgtp



// Seed after: 9947113201368221206,3128299129089410139
