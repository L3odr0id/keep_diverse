// Seed: 12506491258351115114,3128299129089410139

module lssmbw
  (output time kayer [4:1], output reg [0:1][0:3]  qjaxzsk);
  
  
  or bimhh(povlikwrdl, ewergtnunm, qjaxzsk);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:1][0:3]  qjaxzsk -> logic qjaxzsk
  
  
  // Single-driven assigns
  assign kayer = kayer;
  assign qjaxzsk = '{'{'bzz,'b1000,'bx0x,'bz11},'{'bxz11,'b11,'b11z,'b1}};
  
  // Multi-driven assigns
endmodule: lssmbw

module refe
  (output supply0 logic [4:0][1:3][2:0] awo [2:1][1:4], output trireg logic [2:0]  glq);
  
  time otg [4:1];
  
  and jdif(ppkok, ylylhxsej, glq);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   trireg logic [2:0]  glq -> logic glq
  
  lssmbw aighdc(.kayer(otg), .qjaxzsk(vrcwyqnh));
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:1][0:3]  qjaxzsk -> wire logic vrcwyqnh
  
  not soxscnmte(glq, ppkok);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic glq -> trireg logic [2:0]  glq
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign awo = awo;
  assign ppkok = glq;
endmodule: refe

module vup
  ( output logic [1:4][1:0][3:0][3:3]  bpikmojhdo
  , output real keirbad [4:2]
  , input logic [1:2]  rdxmqp
  , input trior logic [4:3][2:3] zchya [1:3]
  , input wand logic [3:4][3:4] szwrue [3:3][4:1]
  );
  
  
  nand raanjrf(cfznmdmjst, mv, pngfwur);
  
  xor upfl(bpikmojhdo, pngfwur, edkzzxlf);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  //   logic bpikmojhdo -> logic [1:4][1:0][3:0][3:3]  bpikmojhdo
  
  not akud(edkzzxlf, mj);
  
  not memmdzvhg(edkzzxlf, mv);
  
  
  // Single-driven assigns
  assign keirbad = '{'b1xx,'bz,'bxx};
  
  // Multi-driven assigns
  assign mv = mj;
endmodule: vup

module boc
  (output supply1 logic [3:4][3:4][1:0][1:0] vm [2:2], input realtime dnr [1:3][3:0], input logic tjhqj);
  
  real eowizjloaj [4:2];
  wand logic [3:4][3:4] gpoe [3:3][4:1];
  trior logic [4:3][2:3] mz [1:3];
  
  and dxmmugxxqw(mfimia, mfimia, mfimia);
  
  xor fxu(ygeqoranj, tjhqj, mfimia);
  
  vup s(.bpikmojhdo(xdbqbz), .keirbad(eowizjloaj), .rdxmqp(hpt), .zchya(mz), .szwrue(gpoe));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   logic [1:4][1:0][3:0][3:3]  bpikmojhdo -> wire logic xdbqbz
  //
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   wire logic hpt -> logic [1:2]  rdxmqp
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: boc



// Seed after: 16560062601981626402,3128299129089410139
