// Seed: 10303539322999713515,3128299129089410139

module nf
  (output trior logic [4:3][4:0][3:2] m [3:4], input bit kvqiiyizxt [2:4][0:0]);
  
  
  not orcwsspuwh(fnd, oxtea);
  
  not t(ogt, nqkuyzlku);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign m = m;
endmodule: nf

module nxeyegttq
  (output time pz, input shortint lepgqgrtt [2:2], input triand logic [2:4][0:0] t [0:4][3:0][3:0], input reg [4:1]  gtoampqtao);
  
  
  
  // Single-driven assigns
  assign pz = 'bz;
  
  // Multi-driven assigns
  assign t = t;
endmodule: nxeyegttq

module jpw
  ( output logic [0:0][3:0] ynzzf [2:4][4:2]
  , output byte cyuuojmjpn
  , input wand logic [2:2][4:1][0:2][2:2] mza [4:2][1:3]
  , input supply1 logic [2:3][4:1][0:0]  mndv
  , input triand logic [2:2][2:1] rps [3:4][3:1][0:2][3:3]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign mndv = '{'{'{'bz},'{'bz1},'{'bxxx1},'{'bxz}},'{'{'b001},'{'bxzx},'{'bzz},'{'bz11}}};
  assign rps = rps;
  assign mza = mza;
endmodule: jpw

module sq
  (output wire logic [0:3][2:3]  wsbeuc);
  
  logic [0:0][3:0] lh [2:4][4:2];
  logic [0:0][3:0] ltmqm [2:4][4:2];
  triand logic [2:2][2:1] owzlclhh [3:4][3:1][0:2][3:3];
  wand logic [2:2][4:1][0:2][2:2] xqridasufn [4:2][1:3];
  triand logic [2:2][2:1] sexknwcmwx [3:4][3:1][0:2][3:3];
  wand logic [2:2][4:1][0:2][2:2] rdifb [4:2][1:3];
  
  jpw ppck(.ynzzf(ltmqm), .cyuuojmjpn(wsbeuc), .mza(rdifb), .mndv(wsbeuc), .rps(sexknwcmwx));
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte cyuuojmjpn -> wire logic [0:3][2:3]  wsbeuc
  
  jpw gzqil(.ynzzf(lh), .cyuuojmjpn(wyiqnmnil), .mza(xqridasufn), .mndv(nhfxs), .rps(owzlclhh));
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte cyuuojmjpn -> wire logic wyiqnmnil
  //
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   wire logic nhfxs -> supply1 logic [2:3][4:1][0:0]  mndv
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nhfxs = wsbeuc;
  assign wyiqnmnil = wsbeuc;
  assign rdifb = rdifb;
endmodule: sq



// Seed after: 13966551278677208945,3128299129089410139
