// Seed: 4170857698512298811,3128299129089410139

module tlk
  ( output trior logic [4:4][1:2][4:1] mdqqkwyja [0:4][2:0][2:1][4:2]
  , output bit ulw [1:1]
  , output logic [1:0] ksptgnzuez [4:3]
  , output reg [3:2][1:4] dns [0:3]
  , input reg ooqcdiyc [4:2][0:0]
  , input tri0 logic vdlck [1:1][0:2][1:4]
  , input byte zrsfbdv [1:2]
  );
  
  
  and wqdxxk(zgybt, cjcux, xgdr);
  
  not vrcz(wmontdg, wsjf);
  
  
  // Single-driven assigns
  assign ulw = ulw;
  assign dns = '{'{'{'b1x,'b0,'b10z10,'bx01x},'{'b01xx1,'b0x1,'bz0xzz,'b0x1zx}},'{'{'b00zz,'b1,'bz,'bzz0x},'{'bz,'b0x000,'b1,'bx0}},'{'{'bz01,'bz101,'bz1000,'b0},'{'bzxz,'b01,'bz,'bz}},'{'{'bxz0,'b0,'bx0,'bz1101},'{'bx0,'b10,'b01,'b0}}};
  assign ksptgnzuez = '{'{'bxxxz,'bzx0z0},'{'b11zz1,'bz1x1}};
  
  // Multi-driven assigns
  assign mdqqkwyja = mdqqkwyja;
  assign cjcux = cjcux;
endmodule: tlk



// Seed after: 3035589897675090996,3128299129089410139
