// Seed: 2461222892141417034,3128299129089410139

module jbynznsyuk
  (output shortreal wadutz [0:1], input logic znz);
  
  
  not yocblbb(tgzyty, znz);
  
  
  // Single-driven assigns
  assign wadutz = wadutz;
  
  // Multi-driven assigns
  assign tgzyty = 'bx;
endmodule: jbynznsyuk

module msupqmjyk
  ( output logic [4:0][3:0][4:2][0:3]  whmw
  , output bit [0:0][2:2][1:3][4:0]  pojjnypdfi
  , output bit [1:2][4:2]  qzn
  , output logic [3:3][4:3][2:1][0:4]  xgzzwfegz
  , input uwire logic [2:3][2:1][4:4][1:1] xnbhzgujsc [4:2][2:4][1:4][3:1]
  );
  
  
  and t(whmw, whmw, pojjnypdfi);
  // warning: implicit conversion of port connection expands from 1 to 240 bits
  //   logic whmw -> logic [4:0][3:0][4:2][0:3]  whmw
  //
  // warning: implicit conversion of port connection truncates from 240 to 1 bits
  //   logic [4:0][3:0][4:2][0:3]  whmw -> logic whmw
  //
  // warning: implicit conversion of port connection truncates from 15 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][2:2][1:3][4:0]  pojjnypdfi -> logic pojjnypdfi
  
  not pvmxoxsej(ibwyphwzpv, gubfkn);
  
  
  // Single-driven assigns
  assign pojjnypdfi = '{'{'{'{'b010,'b1111,'b101,'b011,'b0},'{'b111,'b01,'b00,'b0,'b10},'{'b11010,'b01,'b011,'b101,'b0}}}};
  assign xgzzwfegz = ibwyphwzpv;
  assign qzn = '{'{'b00,'b1010,'b0},'{'b1,'b0111,'b01001}};
  
  // Multi-driven assigns
  assign gubfkn = 'b10;
  assign ibwyphwzpv = 'b1z0x;
endmodule: msupqmjyk



// Seed after: 15147781474257349742,3128299129089410139
