// Seed: 7958188861447328083,3128299129089410139

module imzjv
  (output shortreal xqg [1:2]);
  
  
  not kchdfpycer(tt, oqv);
  
  nand jotzcmwh(tt, qqqwfbbcu, gzo);
  
  not mof(uv, ba);
  
  nand aphhehct(oqv, eqybt, kejj);
  
  
  // Single-driven assigns
  assign xqg = '{'b1,'b1};
  
  // Multi-driven assigns
  assign eqybt = 'bx0x1;
  assign gzo = 'bzz000;
  assign tt = ba;
  assign ba = 'b0;
endmodule: imzjv

module w
  ( output wand logic [4:2] e [3:2]
  , output bit [2:3][3:3][3:4] wlqdil [1:3]
  , output trior logic [1:2][1:3][1:1][4:0] m [4:4][3:3][1:4]
  , input logic [2:1]  l
  , input bit [3:1][3:1][2:2]  axju
  , input bit gbenl
  , input tri logic [2:3][0:4] aonwd [1:1][1:3][3:2][4:0]
  );
  
  shortreal viejto [1:2];
  
  not vzkdevmoqw(b, l);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [2:1]  l -> logic l
  
  not wyuqhgyuw(gaufksvn, axju);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:1][3:1][2:2]  axju -> logic axju
  
  imzjv aw(.xqg(viejto));
  
  
  // Single-driven assigns
  assign wlqdil = wlqdil;
  
  // Multi-driven assigns
  assign e = '{'{'bx1,'bx1,'b0xx1z},'{'b1z1,'bxx0z,'b11z11}};
  assign gaufksvn = 'bx111z;
  assign b = gaufksvn;
  assign aonwd = aonwd;
  assign m = m;
endmodule: w



// Seed after: 13809556470856728717,3128299129089410139
