// Seed: 17120606345259600647,3128299129089410139

module xejv
  ( output wor logic [0:0][0:4][2:3][2:1]  oylynueey
  , output logic [1:3][0:4]  eq
  , output integer e
  , output logic fxuulllgi
  , input bit [0:0][4:0][0:0]  xtpvcd
  );
  
  
  nand us(ex, xtpvcd, dddq);
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][4:0][0:0]  xtpvcd -> logic xtpvcd
  
  not hvqn(reirqbeuq, lkqttegw);
  
  
  // Single-driven assigns
  assign fxuulllgi = eq;
  assign e = 'bz0x0;
  assign eq = oylynueey;
  
  // Multi-driven assigns
  assign oylynueey = '{'{'{'{'b1,'b001},'{'b0,'bz1}},'{'{'bx0,'bx10z1},'{'bz1z,'b1zz0}},'{'{'bz0x,'b0},'{'b0xx1,'bx}},'{'{'b1z1x,'b1z},'{'bz,'bxz}},'{'{'b0,'b1},'{'bz,'b1xzz0}}}};
  assign reirqbeuq = dddq;
  assign ex = lkqttegw;
  assign lkqttegw = oylynueey;
  assign dddq = xtpvcd;
endmodule: xejv



// Seed after: 5762705560976339521,3128299129089410139
