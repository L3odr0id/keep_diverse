// Seed: 10931487316550548278,3128299129089410139

module ufnqkq
  ( output shortreal hqxfhmoae [3:3][0:1]
  , output wor logic [3:4][2:2][0:3]  aztrdcavk
  , input wor logic [4:1][0:4][0:1][4:1] jz [4:0]
  , input uwire logic [3:2][4:2][4:0]  yztybooom
  , input logic [1:1]  t
  );
  
  
  or gcaal(qqslzijnl, t, uo);
  
  or fyy(rj, aztrdcavk, aztrdcavk);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   wor logic [3:4][2:2][0:3]  aztrdcavk -> logic aztrdcavk
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   wor logic [3:4][2:2][0:3]  aztrdcavk -> logic aztrdcavk
  
  xor quojlggxrs(bxmalt, mapliqasi, mapliqasi);
  
  nand bork(aztrdcavk, sciaow, brglxhpvw);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   logic aztrdcavk -> wor logic [3:4][2:2][0:3]  aztrdcavk
  
  
  // Single-driven assigns
  assign hqxfhmoae = hqxfhmoae;
  
  // Multi-driven assigns
  assign bxmalt = aztrdcavk;
  assign aztrdcavk = qqslzijnl;
  assign brglxhpvw = 'b0x1;
  assign rj = bxmalt;
endmodule: ufnqkq

module nzylbwxx
  ( output wire logic [3:1] wzor [0:0][0:0]
  , output trireg logic icxkgmayyp
  , output logic [2:2][3:2][0:0]  rpwgov
  , output triand logic gykozhq
  , input triand logic [2:4][3:1][1:4][2:0] xbk [2:1]
  , input byte piw [0:3][2:0]
  , input supply0 logic [0:2][2:4][2:2][4:2] uyzq [4:4][2:4]
  , input tri0 logic [4:3][1:2] igzc [3:1][4:0][0:3]
  );
  
  
  or b(icxkgmayyp, bqyfkg, fpjoffaan);
  
  and bgvwxcch(rpwgov, icxkgmayyp, t);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic rpwgov -> logic [2:2][3:2][0:0]  rpwgov
  
  and qslcbjfgb(fpjoffaan, rxwrz, hhuidg);
  
  and hjgovos(hllpm, gykozhq, qm);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rxwrz = rxwrz;
  assign hllpm = qm;
  assign icxkgmayyp = 'bz;
  assign bqyfkg = bqyfkg;
endmodule: nzylbwxx



// Seed after: 5862994285518638669,3128299129089410139
