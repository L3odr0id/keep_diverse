// Seed: 13278935458753096407,3128299129089410139

module kliklnrmvx
  ( output wand logic [0:2][0:4][3:0] zellshxjow [1:3]
  , output trior logic [4:4] ftbjmyfrsw [0:3][1:2][0:3][3:2]
  , output logic bvlhjpi
  , input logic [0:4]  gqmhnay
  , input logic t [4:3]
  , input wand logic [2:2][1:4][0:1] thebgzggvc [2:1]
  , input trior logic [2:4][2:4] c [3:4][3:0][4:3]
  );
  
  
  xor gecc(bvlhjpi, bvlhjpi, bvlhjpi);
  
  not va(nbgjtwuk, z);
  
  not lqtu(ttkrqzmcd, tbndinflx);
  
  not ufw(z, bvlhjpi);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: kliklnrmvx

module ady
  ( output reg [1:2]  x
  , output longint ikql
  , input uwire logic [2:2] f [3:0][4:2]
  , input bit [0:3][3:0]  sloxhv
  , input tri logic l
  , input reg [1:1][1:1][4:1]  uqylrzg
  );
  
  
  not hxln(cluy, sloxhv);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:3][3:0]  sloxhv -> logic sloxhv
  
  not qcvbpem(en, uqylrzg);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   reg [1:1][1:1][4:1]  uqylrzg -> logic uqylrzg
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign cluy = 'bz;
  assign en = 'bxz1;
endmodule: ady

module gy
  (input triand logic [1:3][3:1][3:0][0:1] fu [0:2][0:0], input tri0 logic jfh [1:1], input supply0 logic [0:2]  xjumoa);
  
  uwire logic [2:2] mpnikbh [3:0][4:2];
  
  ady lcuqqzra(.x(xjumoa), .ikql(aeezvqu), .f(mpnikbh), .sloxhv(xjumoa), .l(xjumoa), .uqylrzg(xjumoa));
  // warning: implicit conversion of port connection expands from 2 to 3 bits
  //   reg [1:2]  x -> supply0 logic [0:2]  xjumoa
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ikql -> wire logic aeezvqu
  //
  // warning: implicit conversion of port connection expands from 3 to 16 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   supply0 logic [0:2]  xjumoa -> bit [0:3][3:0]  sloxhv
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   supply0 logic [0:2]  xjumoa -> tri logic l
  //
  // warning: implicit conversion of port connection expands from 3 to 4 bits
  //   supply0 logic [0:2]  xjumoa -> reg [1:1][1:1][4:1]  uqylrzg
  
  not s(otrtqudzn, xjumoa);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   supply0 logic [0:2]  xjumoa -> logic xjumoa
  
  or spzt(xjumoa, lwzvhp, lwzvhp);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic xjumoa -> supply0 logic [0:2]  xjumoa
  
  
  // Single-driven assigns
  assign mpnikbh = '{'{'{'bzz},'{'b0z11z},'{'b0}},'{'{'b0z},'{'b000},'{'bz}},'{'{'b0zzx},'{'b00zx},'{'bx}},'{'{'b01x0},'{'bx},'{'b0z100}}};
  
  // Multi-driven assigns
  assign lwzvhp = xjumoa;
  assign fu = fu;
  assign xjumoa = '{'bz,'bx0,'b1};
  assign jfh = jfh;
endmodule: gy

module dsomv
  ( output reg n [2:4]
  , output bit [1:2]  geaoct
  , input supply0 logic [1:3][2:2][4:2] uaitsfej [1:0][3:4]
  , input reg y [2:4]
  , input triand logic jxmltnpnpk [4:0]
  , input reg ol
  );
  
  uwire logic [2:2] guyvvhy [3:0][4:2];
  tri0 logic el [1:1];
  triand logic [1:3][3:1][3:0][0:1] jquxn [0:2][0:0];
  
  nand keul(xiinbdiwc, chibbcwr, chibbcwr);
  
  gy trqzigd(.fu(jquxn), .jfh(el), .xjumoa(geaoct));
  // warning: implicit conversion of port connection expands from 2 to 3 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:2]  geaoct -> supply0 logic [0:2]  xjumoa
  
  ady mjtkhassmb(.x(geaoct), .ikql(ypmf), .f(guyvvhy), .sloxhv(lchfkt), .l(jmospkm), .uqylrzg(xiinbdiwc));
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   reg [1:2]  x -> bit [1:2]  geaoct
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ikql -> wire logic ypmf
  //
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic lchfkt -> bit [0:3][3:0]  sloxhv
  //
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   wire logic xiinbdiwc -> reg [1:1][1:1][4:1]  uqylrzg
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign chibbcwr = geaoct;
  assign el = el;
  assign jquxn = jquxn;
  assign uaitsfej = uaitsfej;
endmodule: dsomv



// Seed after: 14390351302887849332,3128299129089410139
