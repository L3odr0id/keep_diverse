// Seed: 16247055769448328577,3128299129089410139

module fmyedeuj
  ( output trior logic [2:4][0:0][3:2][1:4] okgq [3:2][3:3]
  , output wire logic [4:1][0:3][0:0] ibrb [4:2][4:4]
  , output wand logic [4:4] pryak [1:3][1:0][4:4]
  , input logic [1:2]  yp
  , input logic [2:0][0:0]  ungaf
  , input supply1 logic [4:4] uojkiad [0:3][3:3][3:2]
  );
  
  
  nand skarvuo(oi, s, s);
  
  not f(s, s);
  
  nand mntrcqo(haajzm, q, s);
  
  xor kdxg(zlchjlyszr, camdfbctsd, pmlfhmywuk);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign okgq = okgq;
  assign zlchjlyszr = q;
  assign ibrb = ibrb;
  assign uojkiad = uojkiad;
endmodule: fmyedeuj

module mltmk
  (input reg vkyvmatnw [2:0], input reg [1:1][2:3][3:1]  ojd, input triand logic mgruhq [2:4]);
  
  
  and knquuildu(kwkolyb, ojd, ikfmtfnnb);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   reg [1:1][2:3][3:1]  ojd -> logic ojd
  
  or jbwbxqca(twnks, g, twnks);
  
  xor tjcl(ikfmtfnnb, ikfmtfnnb, dtv);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ikfmtfnnb = g;
endmodule: mltmk

module g
  (output tri0 logic [0:3][0:4][3:3]  euqgkjmiko, input logic [1:3][1:1] ilt [4:2]);
  
  
  and lcvhtb(euqgkjmiko, euqgkjmiko, euqgkjmiko);
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  //   logic euqgkjmiko -> tri0 logic [0:3][0:4][3:3]  euqgkjmiko
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   tri0 logic [0:3][0:4][3:3]  euqgkjmiko -> logic euqgkjmiko
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   tri0 logic [0:3][0:4][3:3]  euqgkjmiko -> logic euqgkjmiko
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: g



// Seed after: 4730330285713594232,3128299129089410139
