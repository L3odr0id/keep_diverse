// Seed: 3118380402852848225,3128299129089410139

module epsbfthuq
  (output logic [3:1][1:2]  okiumnjw, output bit tuafcrfqgo, output trior logic [1:2] btmiwshot [3:1][4:4][3:1][3:4]);
  
  
  not rgx(pdmtxt, gxzndoeil);
  
  or chhls(tuafcrfqgo, ferkwhus, gxzndoeil);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic tuafcrfqgo -> bit tuafcrfqgo
  
  
  // Single-driven assigns
  assign okiumnjw = okiumnjw;
  
  // Multi-driven assigns
  assign btmiwshot = btmiwshot;
endmodule: epsbfthuq



// Seed after: 1276793512140722276,3128299129089410139
