// Seed: 8441463012171610221,3128299129089410139

module fkng
  ( output tri0 logic [1:0][1:0] tcpb [3:1][2:2][0:4]
  , output int mgjycuwj [4:2]
  , input bit [1:0] q [2:3]
  , input tri1 logic [3:2] emfah [1:2][1:0][1:2]
  , input supply1 logic [3:2][0:1][3:4][3:4] vh [3:4]
  , input real xjh [0:0]
  );
  
  
  and ucblnhpasc(dvmctbe, azsws, azsws);
  
  or lmrtz(py, qckdtnyk, keej);
  
  not f(dvmctbe, azsws);
  
  xor ytqj(kettayvd, dvmctbe, ttw);
  
  
  // Single-driven assigns
  assign mgjycuwj = '{'b100,'b0000,'b101};
  
  // Multi-driven assigns
  assign tcpb = tcpb;
  assign dvmctbe = 'b0;
  assign ttw = azsws;
  assign azsws = ttw;
  assign py = azsws;
endmodule: fkng

module xadvv
  ( output reg [0:2][1:1]  ckt
  , input tri0 logic czfmqebhn [0:0]
  , input bit [3:1][0:2]  m
  , input triand logic [0:4][3:0][1:2][2:1] wy [0:0][2:3][0:2]
  , input tri logic [2:0] zboxxis [0:4][1:2][4:1][3:3]
  );
  
  
  not tsseff(ckt, ckt);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic ckt -> reg [0:2][1:1]  ckt
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][1:1]  ckt -> logic ckt
  
  not zpljgix(iknoqsqgfm, mwokb);
  
  not ojglusbiqw(lklxo, ckt);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][1:1]  ckt -> logic ckt
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: xadvv



// Seed after: 6882737065302465407,3128299129089410139
