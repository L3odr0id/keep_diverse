// Seed: 6882737065302465407,3128299129089410139

module gvbnbvvrfw
  ( output uwire logic [4:4][0:0] yrrshvik [0:0]
  , output bit [0:3][1:0][1:3] wrxfoufw [4:4]
  , output tri1 logic [2:2]  ipqffsdnxk
  , output int sopczjg
  , input uwire logic [3:0][3:4] zekgn [3:1][3:3]
  , input logic [3:0]  jtqlupj
  );
  
  
  not yr(djzfqxcjj, ykwpppsgb);
  
  not rq(b, qwu);
  
  or hgyvup(djzfqxcjj, ipqffsdnxk, ykwpppsgb);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: gvbnbvvrfw



// Seed after: 10573157214128529296,3128299129089410139
