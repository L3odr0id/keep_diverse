// Seed: 1536635323995096370,3128299129089410139

module iynxjytram
  (output shortint dxgtc);
  
  
  not jssegzpbup(dxgtc, dxgtc);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic dxgtc -> shortint dxgtc
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint dxgtc -> logic dxgtc
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: iynxjytram

module rufxlngeye
  ( output triand logic [3:0][0:3] ylp [3:3][3:0][1:1][0:1]
  , output tri logic [4:4][3:3][4:3][4:3] ovqyhzl [3:3]
  , input bit [1:3][1:3][3:2][0:1]  vh
  , input tri1 logic [1:1][2:3][2:2] ttnmeikzcf [3:0][1:0][1:3]
  , input time u [3:3]
  , input real lujc
  );
  
  
  not gffazco(r, lujc);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real lujc -> logic lujc
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ovqyhzl = ovqyhzl;
  assign r = 'bxx0xx;
  assign ttnmeikzcf = ttnmeikzcf;
  assign ylp = ylp;
endmodule: rufxlngeye



// Seed after: 430576150281111274,3128299129089410139
