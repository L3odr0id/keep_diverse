// Seed: 2428324134062495893,3128299129089410139

module vk
  (output bit [4:1][1:1][2:2][1:4]  cwx, output shortreal gey [0:0][1:2], input wire logic [1:0][2:2][4:1] tikr [2:2][4:2][0:1][2:2]);
  
  
  not hhugvquhv(cwx, jotvqzmqs);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic cwx -> bit [4:1][1:1][2:2][1:4]  cwx
  
  not dosvqanbs(jotvqzmqs, tnngpi);
  
  
  // Single-driven assigns
  assign gey = gey;
  
  // Multi-driven assigns
  assign tnngpi = cwx;
  assign tikr = tikr;
endmodule: vk



// Seed after: 17774132640328010878,3128299129089410139
