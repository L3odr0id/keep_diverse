// Seed: 11532771568697646238,3128299129089410139

module m
  ( output tri0 logic [0:2][3:2][0:3][0:2] li [3:0][1:4][1:2][2:1]
  , output bit mwwn [1:2]
  , input logic ccyegpbg [2:0]
  , input uwire logic [1:3][2:1][3:2][4:2] z [4:4][4:4][3:3]
  , input tri0 logic dgm [0:4][3:1]
  , input triand logic [4:0][1:0][1:2][4:4] qa [0:0][4:2][0:2]
  );
  
  
  not ebsqw(zxbzf, zxbzf);
  
  not hqijqwc(jy, jy);
  
  nand hhsepxvv(jy, kroeyjnbnc, ovsmlmufum);
  
  xor dlnwxu(csoct, zxbzf, zxbzf);
  
  
  // Single-driven assigns
  assign mwwn = mwwn;
  
  // Multi-driven assigns
  assign li = li;
  assign zxbzf = 'bx011x;
endmodule: m

module prmymrhi
  ( output wor logic [0:4][3:1] mwxfmqmk [1:2][1:1][2:4][3:0]
  , output logic [4:4][0:1][4:2][1:4]  rbsi
  , output integer zpadxjvq
  , input logic [3:0]  ilwqym
  , input tri logic [1:4][2:4] auramgbmnb [3:1]
  , input wire logic [2:0][1:2][0:1] nftyyzhx [4:1][4:1][0:4][3:1]
  );
  
  
  
  // Single-driven assigns
  assign rbsi = '{'{'{'{'b0,'bx,'b1,'b1x1},'{'b1,'bx1x0,'bz,'bz},'{'b0x,'b10,'bx0xxz,'bx0xz}},'{'{'bx1,'bxzzx1,'b0110,'b0zz1},'{'bz1,'b1x0zz,'b1z,'b1xxx1},'{'b0zxzz,'bx11,'bx11,'bzz101}}}};
  
  // Multi-driven assigns
  assign mwxfmqmk = mwxfmqmk;
  assign nftyyzhx = nftyyzhx;
  assign auramgbmnb = '{'{'{'bx1xxx,'bz1z,'b0},'{'bzz0x,'bz0z1,'b0},'{'bz00,'bx01,'bxx11z},'{'bz01zz,'b00z,'b1z0}},'{'{'b00zx,'bxxxx,'b1z},'{'b0x,'bx0z0,'bz0},'{'bxzzz,'b11zz,'b11x1},'{'b0,'bzx1zz,'b0}},'{'{'bx1,'b1,'bx0},'{'bzxx0,'b011x,'b111x},'{'b000xz,'b10,'bxzxz},'{'bzz0z0,'bx0xxx,'b0zz1x}}};
endmodule: prmymrhi

module sqjlrl
  (output tri logic [0:2][4:2][3:4]  qt, input bit [3:1]  jbkiyshric, input wand logic [2:3][0:4] rsrfyjble [2:2][2:3][2:4]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign qt = qt;
  assign rsrfyjble = rsrfyjble;
endmodule: sqjlrl



// Seed after: 5893021453546226726,3128299129089410139
