// Seed: 7084504391126471160,3128299129089410139

module eyk
  (output triand logic [1:1][2:3]  fcu, input supply0 logic [4:0]  oqzmoesoqo);
  
  
  nand rzjtmlfpri(fcu, w, w);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic fcu -> triand logic [1:1][2:3]  fcu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign oqzmoesoqo = '{'bz1,'b1,'b1zx,'bx,'b0};
  assign w = 'bzzx10;
  assign fcu = fcu;
endmodule: eyk

module mkjozxh
  ( output reg [3:1][4:3]  jxdnjza
  , output uwire logic aveyi [4:0][2:3][3:0]
  , output logic [0:4][1:3]  lpmezxeho
  , output reg [1:1] d [0:1]
  , input trireg logic [0:3][0:0][0:4] ye [3:2][2:3][3:4]
  , input tri logic [4:2][2:4] wsnokqlm [2:2][2:2][1:3]
  );
  
  
  nand aogp(joacltk, joacltk, jxdnjza);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   reg [3:1][4:3]  jxdnjza -> logic jxdnjza
  
  or f(x, xyzd, jxdnjza);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   reg [3:1][4:3]  jxdnjza -> logic jxdnjza
  
  nand mo(wunsagt, lpmezxeho, dh);
  // warning: implicit conversion of port connection truncates from 15 to 1 bits
  //   logic [0:4][1:3]  lpmezxeho -> logic lpmezxeho
  
  not pscylwwcg(kro, xyzd);
  
  
  // Single-driven assigns
  assign jxdnjza = joacltk;
  assign lpmezxeho = '{'{'bz0111,'bz00xx,'b011},'{'bx,'bzx,'b1x101},'{'b01,'bzz,'b111},'{'bx0zzx,'b1z1,'bz0z},'{'b0,'bz0z0,'b1}};
  assign aveyi = aveyi;
  
  // Multi-driven assigns
  assign ye = ye;
  assign joacltk = 'bx1;
  assign xyzd = 'b0;
endmodule: mkjozxh

module itjd
  ( output reg [4:4]  ab
  , output logic [2:1][3:0][2:1]  xaeximp
  , output tri logic [4:4] xyzbhm [1:2][0:2][1:2][2:0]
  , output logic [1:1][2:2][4:3]  olurwydwvh
  , input tri0 logic [0:1][4:0][0:3][0:4] eursa [1:4]
  , input reg [2:4]  ptatr
  , input logic [4:4][3:3][0:4] tmcntnxmz [2:1]
  , input bit [1:2][0:3]  dowhc
  );
  
  
  or jqyadump(em, xaeximp, ptatr);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   logic [2:1][3:0][2:1]  xaeximp -> logic xaeximp
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [2:4]  ptatr -> logic ptatr
  
  
  // Single-driven assigns
  assign olurwydwvh = ab;
  
  // Multi-driven assigns
endmodule: itjd



// Seed after: 3118380402852848225,3128299129089410139
