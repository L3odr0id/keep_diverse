// Seed: 15147781474257349742,3128299129089410139

module fdnt
  ( output wire logic [1:2] kwcgsfl [0:2]
  , input tri logic [2:0] qftdqraxr [3:2][1:3][4:1][4:4]
  , input supply0 logic it [4:3]
  , input int no
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: fdnt

module pnqzbr
  ( output trireg logic [3:3][2:3][0:0][0:3]  hsjtwdgiir
  , output byte n
  , input tri logic [1:1][1:2][3:3] f [3:2]
  , input integer spuwhyfb
  , input supply0 logic [2:0][3:4] puavwkjuhv [4:0][0:4][0:3]
  );
  
  
  
  // Single-driven assigns
  assign n = spuwhyfb;
  
  // Multi-driven assigns
  assign hsjtwdgiir = hsjtwdgiir;
  assign f = f;
endmodule: pnqzbr



// Seed after: 2428324134062495893,3128299129089410139
