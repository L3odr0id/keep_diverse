// Seed: 6580800625636262848,3128299129089410139

module xyfbg
  (input longint uzmsulku [2:2], input tri1 logic [1:1][4:4][3:4]  vzvpgn, input reg [2:2]  khfbaqoqa);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign vzvpgn = vzvpgn;
endmodule: xyfbg



// Seed after: 4919911431090630944,3128299129089410139
