// Seed: 11334337321803779299,3128299129089410139

module uwlcs
  ( output logic [4:0]  kbwuiwc
  , output bit [4:2][2:4]  byemmnmvtj
  , input tri1 logic osoflydb
  , input shortint g
  , input logic [4:3][2:2][3:2][0:2]  tsmvywyjxp
  );
  
  
  not xgawhdzvq(kbwuiwc, byemmnmvtj);
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   logic kbwuiwc -> logic [4:0]  kbwuiwc
  //
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:2][2:4]  byemmnmvtj -> logic byemmnmvtj
  
  not yqk(hvqxncj, osoflydb);
  
  not jy(byemmnmvtj, gtfjlqebp);
  // warning: implicit conversion of port connection expands from 1 to 9 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic byemmnmvtj -> bit [4:2][2:4]  byemmnmvtj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign osoflydb = kbwuiwc;
  assign hvqxncj = 'b0;
  assign gtfjlqebp = 'b101;
endmodule: uwlcs



// Seed after: 8441463012171610221,3128299129089410139
