// Seed: 3969165351885200449,3128299129089410139

module sootvnwy
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: sootvnwy

module cy
  (output tri0 logic [0:1] algpsbk [4:1], output bit ucdbg, output real uufyoa, input logic [4:3][4:4] foivmo [3:0]);
  
  
  or yoysy(fuztjuvrv, ucdbg, oapffjb);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit ucdbg -> logic ucdbg
  
  sootvnwy lhvfydx();
  
  not naowxhfru(uufyoa, qyvfdmrqib);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic uufyoa -> real uufyoa
  
  
  // Single-driven assigns
  assign ucdbg = 'b01;
  
  // Multi-driven assigns
  assign fuztjuvrv = 'b0z;
  assign oapffjb = 'bx0x;
  assign algpsbk = algpsbk;
endmodule: cy

module dvnrcjn
  (output real lytckhx, output supply0 logic [3:2][3:2][1:0][0:1] ymra [1:3], input reg [1:2]  cjnun);
  
  logic [4:3][4:4] b [3:0];
  
  cy hhby(.algpsbk(b), .ucdbg(grnqhykl), .uufyoa(d), .foivmo(b));
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit ucdbg -> wire logic grnqhykl
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real uufyoa -> wire logic d
  
  
  // Single-driven assigns
  assign lytckhx = 'bx00z;
  
  // Multi-driven assigns
  assign ymra = ymra;
  assign grnqhykl = cjnun;
  assign d = 'b1;
endmodule: dvnrcjn

module usnq
  (output trireg logic [0:4][3:4][4:1][1:0]  dblx, output trireg logic [1:2] ygjvupamjz [3:1][2:4][2:2]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dblx = '{'{'{'{'b1,'b00x0z},'{'b011x,'bz00},'{'bx0z00,'bzxz},'{'b010x0,'bz111}},'{'{'b0,'b0110x},'{'bx,'b11zzx},'{'bx0,'bzxx},'{'bz0x,'bzz11}}},'{'{'{'bz0zx0,'bxx1},'{'b0xxxx,'bzx1},'{'bzzzx,'bx0xx0},'{'b0,'bz1zx}},'{'{'b0zzx,'bx00x},'{'b001zx,'bz0},'{'bx010,'bzxx},'{'b1,'b1}}},'{'{'{'b11,'bz1xzx},'{'bz0x,'bxx},'{'bzz01z,'b1},'{'bx,'bxxx0}},'{'{'bzz00,'bzzx1},'{'bxzx10,'b1z0},'{'b0,'b0x},'{'b0x0,'b0}}},'{'{'{'bx01z,'bzx00},'{'bxxzx,'b0zz},'{'bx0,'b0z0z1},'{'bxz,'b0xzz0}},'{'{'b0z0,'b10zz},'{'bx0xz0,'b10z},'{'bx111,'bx11},'{'bzzz,'b0z010}}},'{'{'{'b0,'b01z0},'{'bzzxxz,'b101},'{'bx1,'bzz10z},'{'b1,'b11xz}},'{'{'bx10xx,'b1},'{'b00,'b1x0},'{'b1,'b00},'{'bx1,'bz01zz}}}};
  assign ygjvupamjz = ygjvupamjz;
endmodule: usnq



// Seed after: 4427233426964322947,3128299129089410139
