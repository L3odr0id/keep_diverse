// Seed: 9058340612855349718,3128299129089410139

module wdxyoedogi
  ( output triand logic [3:3][3:2][4:2] jwuk [3:2][4:1]
  , input bit [2:4][3:4][2:1] ewoacsvxxu [0:3]
  , input uwire logic [2:0][0:0][0:3][2:3] nkhmytgi [4:2]
  , input trireg logic [2:4] nueszgvjlk [4:0]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: wdxyoedogi

module e
  (output uwire logic [0:0][0:4] jzsu [3:3][4:4][1:0][0:4], input supply1 logic ld [3:3]);
  
  
  or uvhvmgri(d, mqm, mqm);
  
  nand lbm(du, mqm, glvrpnctk);
  
  not ookp(saofqmv, d);
  
  
  // Single-driven assigns
  assign jzsu = jzsu;
  
  // Multi-driven assigns
endmodule: e

module yehuw
  ( output tri0 logic tappmu
  , output trior logic jrpj [4:2][3:4][2:4][0:4]
  , output supply1 logic [2:2] us [1:3][0:1]
  , input tri logic [0:0][0:3] nrk [3:0][2:3]
  , input shortreal fgcyi
  , input wor logic [2:2][2:1] hij [3:3][2:4][3:3]
  , input trior logic [4:1][0:0][2:2] oojxjjcxrw [4:0][2:2]
  );
  
  
  nand bonulswq(zceovjw, tappmu, ifgl);
  
  and eovzddysw(tappmu, elegar, qgzuxsik);
  
  not ebwxec(zb, tappmu);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zceovjw = 'b1z;
  assign tappmu = 'bzz;
  assign jrpj = '{'{'{'{'b110xx,'b11,'b001,'bxzz0,'b1zx},'{'bxzz,'bx1zz,'b1xxx,'bz010x,'b1xx},'{'b11,'bz1,'bxzx0,'b0,'b1}},'{'{'bx11,'b00,'bz0xxx,'b1,'b00},'{'b1x,'bx00z1,'bz1xz,'bzz0,'b1z},'{'b0,'b0,'bx,'bz,'bx11z0}}},'{'{'{'bx,'b1z0,'bz1,'bxzxz,'b10x},'{'b1z,'bz1z,'b111x,'b1,'bxz0zz},'{'bx0,'b1x,'b10x0,'bx,'b001}},'{'{'b01zx1,'bzx0,'b1x1,'b0,'bxz00},'{'b0z0x,'b1,'bx001z,'b00x,'bx},'{'b0,'b10,'bx1,'b110zx,'b1}}},'{'{'{'bxz,'b0z,'b100,'b0z01,'bx},'{'b11z,'b00,'bzz0,'bx01z,'bz},'{'b0xz1x,'b1,'bxxzz,'bx0,'bz}},'{'{'bxz1z1,'bx11z,'bxz,'bx,'bxzz},'{'bzz1zx,'bz,'bzxz1z,'bxxxx1,'bzxz},'{'b1z1xz,'bx,'b00x1,'bx1zx,'bz}}}};
  assign qgzuxsik = qgzuxsik;
endmodule: yehuw



// Seed after: 16397190719548895153,3128299129089410139
