// Seed: 18305973876864763085,3128299129089410139

module klksylif
  ( input reg [1:3][0:1]  ngzaw
  , input logic [4:2][4:3][4:4]  gfmocscbux
  , input reg [0:2][3:0] zeruk [1:3]
  , input tri logic [2:0][4:1] hzh [4:2][1:1]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hzh = hzh;
endmodule: klksylif



// Seed after: 13160880725827085634,3128299129089410139
