// Seed: 686311863841549876,3128299129089410139

module vfneom
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: vfneom

module mbgwabqt
  ( output tri1 logic [2:2][1:3][2:2]  qulmwa
  , input supply1 logic [4:3][3:2][3:2] meydx [1:2]
  , input tri0 logic xwccot
  , input bit [2:0][0:2] fr [1:2]
  , input bit [1:3][2:2][4:0]  ydws
  );
  
  
  or ufy(qulmwa, qulmwa, qulmwa);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic qulmwa -> tri1 logic [2:2][1:3][2:2]  qulmwa
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qulmwa
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qulmwa
  
  not zdlcc(ycosloucl, qulmwa);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qulmwa
  
  and akaj(kmah, qulmwa, qulmwa);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qulmwa
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qulmwa
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kmah = 'b0x010;
  assign xwccot = 'bxxzx;
  assign qulmwa = '{'{'{'bx},'{'b00zz},'{'bzx}}};
  assign meydx = meydx;
  assign ycosloucl = qulmwa;
endmodule: mbgwabqt

module qu
  ( output bit cbwi
  , output supply1 logic [2:1][1:4][0:4] jlb [3:3][0:1][4:4]
  , output reg [3:4]  tdcveqn
  , output reg [1:1][4:2][4:3]  fhzxlc
  );
  
  
  not xtbhog(kcnu, tdcveqn);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   reg [3:4]  tdcveqn -> logic tdcveqn
  
  
  // Single-driven assigns
  assign cbwi = 'b00;
  assign fhzxlc = '{'{'{'b0z,'b0x},'{'b11,'bz},'{'b010,'bx0x11}}};
  assign tdcveqn = '{'b0,'bz0};
  
  // Multi-driven assigns
endmodule: qu

module oyuu
  ( output logic qmdqpmrq
  , output realtime hngli [1:3]
  , output tri logic johkojmndw
  , output reg [0:2]  oumjz
  , input int updjipgzv
  , input real sq
  , input tri logic so [0:0][0:0]
  );
  
  bit [2:0][0:2] uuhms [1:2];
  supply1 logic [4:3][3:2][3:2] byaxlpc [1:2];
  
  and vljcuaxkgs(htd, wkdch, qmdqpmrq);
  
  mbgwabqt htgdwngrew(.qulmwa(qmdqpmrq), .meydx(byaxlpc), .xwccot(j), .fr(uuhms), .ydws(hiydbmmd));
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri1 logic [2:2][1:3][2:2]  qulmwa -> logic qmdqpmrq
  //
  // warning: implicit conversion of port connection expands from 1 to 15 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic hiydbmmd -> bit [1:3][2:2][4:0]  ydws
  
  nand zgrbmxurjs(johkojmndw, qmdqpmrq, htd);
  
  vfneom fuqduu();
  
  
  // Single-driven assigns
  assign hngli = hngli;
  assign uuhms = uuhms;
  assign oumjz = qmdqpmrq;
  
  // Multi-driven assigns
  assign johkojmndw = j;
  assign hiydbmmd = 'bz;
endmodule: oyuu



// Seed after: 13299826562397828311,3128299129089410139
