// Seed: 5862994285518638669,3128299129089410139

module ssjftj
  ( output tri1 logic [2:2] il [4:4]
  , input supply0 logic [1:4][2:3] uge [1:4][2:0][4:2][4:0]
  , input wire logic [3:3][4:4][0:3][1:3]  gzefx
  );
  
  
  not l(nsekaylq, gzefx);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   wire logic [3:3][4:4][0:3][1:3]  gzefx -> logic gzefx
  
  and jv(bjzabehpxn, bjzabehpxn, gzefx);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   wire logic [3:3][4:4][0:3][1:3]  gzefx -> logic gzefx
  
  nand levmk(gzefx, hypbr, gzefx);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic gzefx -> wire logic [3:3][4:4][0:3][1:3]  gzefx
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   wire logic [3:3][4:4][0:3][1:3]  gzefx -> logic gzefx
  
  or lkixuertf(gzefx, gzefx, nsekaylq);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic gzefx -> wire logic [3:3][4:4][0:3][1:3]  gzefx
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   wire logic [3:3][4:4][0:3][1:3]  gzefx -> logic gzefx
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign il = il;
  assign gzefx = gzefx;
endmodule: ssjftj

module ienl
  ( output wor logic [3:4][0:2][1:4][1:2] dndnrimj [4:0]
  , output bit [2:1][0:1][4:1]  svqs
  , input uwire logic [0:3][1:1][1:3][2:2] pkamimx [0:4][1:3]
  , input tri logic [2:0][1:4][4:1] ucuirdie [3:2][3:4][0:4]
  , input wand logic [4:4][3:2][2:1] n [3:1]
  , input supply1 logic wlptbgnx [2:1][4:1][2:3]
  );
  
  tri1 logic [2:2] sr [4:4];
  supply0 logic [1:4][2:3] jyasif [1:4][2:0][4:2][4:0];
  
  not onvbdq(fzuwnehio, mruwf);
  
  or klejgvypt(wrfpfhtur, hijcleala, svqs);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1][0:1][4:1]  svqs -> logic svqs
  
  ssjftj gk(.il(sr), .uge(jyasif), .gzefx(uncuvouak));
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic uncuvouak -> wire logic [3:3][4:4][0:3][1:3]  gzefx
  
  or mmo(qc, svqs, aqcyphezk);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1][0:1][4:1]  svqs -> logic svqs
  
  
  // Single-driven assigns
  assign svqs = svqs;
  
  // Multi-driven assigns
  assign ucuirdie = ucuirdie;
  assign dndnrimj = dndnrimj;
  assign n = '{'{'{'{'b001,'bzzz1},'{'bxz0,'bx}}},'{'{'{'bx0zz,'bz1x},'{'b001,'bxxx0}}},'{'{'{'bxxzx1,'b111},'{'b1zz0z,'b1}}}};
  assign sr = '{'{'bx1x}};
  assign mruwf = svqs;
endmodule: ienl



// Seed after: 9407371298728588963,3128299129089410139
