// Seed: 9741254061059762472,3128299129089410139

module lrlnswuh
  ( output bit [3:1][3:1]  lqcggv
  , output uwire logic [3:0][3:3] zjq [4:2][0:0][4:4]
  , input triand logic ynt [3:1][4:0][0:0][4:4]
  , input supply0 logic [3:2][4:2][2:1][4:0] ltgs [1:1][1:3][0:4]
  );
  
  
  not s(vigcqlozod, birgfc);
  
  xor mnjslfzvty(ldmefm, lqcggv, vpeqozlbai);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:1][3:1]  lqcggv -> logic lqcggv
  
  or bz(n, lqcggv, vpeqozlbai);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:1][3:1]  lqcggv -> logic lqcggv
  
  xor tsbl(lqcggv, lqcggv, vpeqozlbai);
  // warning: implicit conversion of port connection expands from 1 to 9 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic lqcggv -> bit [3:1][3:1]  lqcggv
  //
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:1][3:1]  lqcggv -> logic lqcggv
  
  
  // Single-driven assigns
  assign zjq = zjq;
  
  // Multi-driven assigns
  assign ltgs = ltgs;
  assign ynt = '{'{'{'{'b01}},'{'{'bxxz01}},'{'{'b0010}},'{'{'bxx}},'{'{'b101zx}}},'{'{'{'bzxxx1}},'{'{'b11}},'{'{'b1}},'{'{'bx}},'{'{'bxz}}},'{'{'{'b1zzz}},'{'{'b1xx}},'{'{'bzx0}},'{'{'bzx0}},'{'{'bz}}}};
  assign birgfc = 'bxx0;
  assign vpeqozlbai = 'b0;
  assign n = 'b01x01;
endmodule: lrlnswuh

module jrdmktnn
  (input wor logic [4:2]  shvovwrd, input int puuxrcto, input longint luf);
  
  
  xor isgaw(shvovwrd, shvovwrd, puuxrcto);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic shvovwrd -> wor logic [4:2]  shvovwrd
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wor logic [4:2]  shvovwrd -> logic shvovwrd
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int puuxrcto -> logic puuxrcto
  
  nand muwaugkm(shvovwrd, luf, luf);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic shvovwrd -> wor logic [4:2]  shvovwrd
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint luf -> logic luf
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint luf -> logic luf
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign shvovwrd = '{'b1,'b01x,'bzxx};
endmodule: jrdmktnn

module eq
  ( output int tm [2:3][4:4]
  , output wire logic [3:1] vmhequkl [3:1][3:1][1:0]
  , output tri logic [1:0][1:4][2:1] mcylcuw [2:0][3:4][1:1][4:3]
  );
  
  
  xor ngl(mwjaa, td, td);
  
  not zfboqxzt(aiucnf, ucvvj);
  
  
  // Single-driven assigns
  assign tm = tm;
  
  // Multi-driven assigns
endmodule: eq



// Seed after: 4170857698512298811,3128299129089410139
