// Seed: 10573157214128529296,3128299129089410139

module h
  ( output uwire logic [3:0][2:3][3:0][1:4]  qziljglti
  , output trior logic [3:4][1:3][3:4] okitugarik [4:1][1:0][3:2][3:1]
  , output bit [0:3]  glqytyaeeb
  , input logic [0:0][2:0] pdkeknp [0:2]
  , input trireg logic [1:1][2:2][0:0] gnm [2:4][3:0]
  , input wand logic [2:3][4:2][4:1][1:4]  xekagvkf
  , input trireg logic [0:2][0:3] e [0:2][1:4][2:4][2:1]
  );
  
  
  xor wufaeeerr(jgsipuow, m, glqytyaeeb);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:3]  glqytyaeeb -> logic glqytyaeeb
  
  nand eqy(t, ywhcvlvsc, gjei);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign e = e;
  assign gnm = gnm;
  assign t = glqytyaeeb;
endmodule: h

module mwmnifa
  ();
  
  
  nand ho(cumdprt, j, cumdprt);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: mwmnifa



// Seed after: 686311863841549876,3128299129089410139
