// Seed: 17774132640328010878,3128299129089410139

module pln
  ( output logic [2:0][3:3][4:3] ueunlqiosb [2:1]
  , output real b
  , output uwire logic [0:3][3:2][2:2][0:4] iemg [2:1][3:4][4:3][1:3]
  , output bit [0:3][4:4] da [2:1]
  , input logic [2:2][2:4] kmaetucw [4:3]
  );
  
  
  and udijxugj(rt, b, b);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real b -> logic b
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real b -> logic b
  
  xor eih(xtxsrveekf, rt, xtxsrveekf);
  
  
  // Single-driven assigns
  assign ueunlqiosb = '{'{'{'{'bzx,'bz}},'{'{'bxzz0,'bzz1}},'{'{'b0,'b10z}}},'{'{'{'bz010z,'bx0x1}},'{'{'bzxxx0,'bxz}},'{'{'bx1x0x,'b1z0}}}};
  assign b = 'b1zz0;
  assign da = '{'{'{'b00111},'{'b000},'{'b10},'{'b11110}},'{'{'b10101},'{'b001},'{'b00},'{'b1}}};
  
  // Multi-driven assigns
  assign rt = 'bx0zz;
  assign xtxsrveekf = xtxsrveekf;
endmodule: pln

module mdr
  ( output reg [3:1][3:3][3:2][1:0]  ynxq
  , output tri logic [2:2][4:3] j [2:3][2:4][4:1][4:0]
  , input tri1 logic [3:4][3:0] hkr [2:0][4:0]
  , input logic [2:0][1:1][4:2]  tjflm
  , input logic htphgbjkr [1:4]
  );
  
  bit [0:3][4:4] m [2:1];
  uwire logic [0:3][3:2][2:2][0:4] mg [2:1][3:4][4:3][1:3];
  logic [2:0][3:3][4:3] w [2:1];
  logic [2:2][2:4] eoec [4:3];
  
  or wp(mfpmrpx, ab, mfpmrpx);
  
  pln eees(.ueunlqiosb(w), .b(ynxq), .iemg(mg), .da(m), .kmaetucw(eoec));
  // warning: implicit conversion of port connection truncates from 64 to 12 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real b -> reg [3:1][3:3][3:2][1:0]  ynxq
  
  nand cw(wsehbcoz, ynxq, ynxq);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [3:1][3:3][3:2][1:0]  ynxq -> logic ynxq
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [3:1][3:3][3:2][1:0]  ynxq -> logic ynxq
  
  and swf(ab, hltjiemvoi, tjflm);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  //   logic [2:0][1:1][4:2]  tjflm -> logic tjflm
  
  
  // Single-driven assigns
  assign eoec = eoec;
  
  // Multi-driven assigns
  assign j = j;
  assign ab = tjflm;
endmodule: mdr



// Seed after: 8699459758548135104,3128299129089410139
