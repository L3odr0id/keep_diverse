// Seed: 574283273884231197,3128299129089410139

module imadsbksr
  ( output triand logic [0:3] flfdgehflp [2:2][4:1][0:2][4:4]
  , output bit [4:0][1:0] jqrqpsgqnh [4:0]
  , input reg de
  , input triand logic [0:4][4:4][4:2] dvglr [2:0]
  , input supply1 logic [2:2][0:0]  zn
  );
  
  
  not w(gorrpcvp, zn);
  
  
  // Single-driven assigns
  assign jqrqpsgqnh = '{'{'{'b01,'b1},'{'b1010,'b1010},'{'b0110,'b1},'{'b001,'b01001},'{'b00,'b0000}},'{'{'b01,'b11000},'{'b000,'b110},'{'b10111,'b100},'{'b00011,'b11010},'{'b111,'b0}},'{'{'b0,'b1},'{'b10,'b0100},'{'b10100,'b1},'{'b0,'b0000},'{'b01010,'b0}},'{'{'b110,'b010},'{'b01010,'b01},'{'b100,'b1011},'{'b100,'b01011},'{'b11111,'b01}},'{'{'b10010,'b0},'{'b0,'b01010},'{'b00110,'b10},'{'b01,'b1},'{'b1100,'b11}}};
  
  // Multi-driven assigns
  assign dvglr = '{'{'{'{'b1x1,'bxzx01,'bz011x}},'{'{'b0zz,'bx1zxz,'b1x}},'{'{'b0,'b00z01,'b111xz}},'{'{'bz0,'bxz0,'b0zxx}},'{'{'bx1z,'bxxzx,'bz1zz}}},'{'{'{'b1,'b1,'b0x10x}},'{'{'bx0z0x,'bz01x,'b01}},'{'{'b1,'b0,'bzxz01}},'{'{'bx0,'b110,'b01}},'{'{'b1xx,'b1xzz1,'bz00xx}}},'{'{'{'b0,'bx1,'bzz1}},'{'{'bx0,'bz01,'b11z1}},'{'{'bxxx,'bz,'b1z0z1}},'{'{'b101xx,'bx,'b010}},'{'{'b011z1,'b100x,'b1x}}}};
  assign flfdgehflp = flfdgehflp;
  assign zn = '{'{'b11z}};
endmodule: imadsbksr

module w
  ( output uwire logic [4:2][0:2] xpb [1:3][1:0][4:2][0:2]
  , input tri1 logic [3:1][0:2][0:4][1:2]  rqlxilvgw
  , input integer zxh
  , input supply1 logic [3:4][0:2][2:1][0:3] fgsbjey [1:1]
  , input longint qox
  );
  
  
  not s(rqlxilvgw, zxh);
  // warning: implicit conversion of port connection expands from 1 to 90 bits
  //   logic rqlxilvgw -> tri1 logic [3:1][0:2][0:4][1:2]  rqlxilvgw
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer zxh -> logic zxh
  
  
  // Single-driven assigns
  assign xpb = xpb;
  
  // Multi-driven assigns
endmodule: w



// Seed after: 5290427713959618967,3128299129089410139
