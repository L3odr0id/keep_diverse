// Seed: 4868562018233217693,3128299129089410139

module lgogd
  ( output logic [1:1][4:3]  wgaioirl
  , input logic ur [2:4]
  , input trireg logic [2:0][4:2][4:4] ercrh [2:4][3:0][1:3]
  , input tri logic [2:2][0:0]  gbpuekkj
  , input supply1 logic [0:3][2:2][3:4] ceegabuwg [4:2]
  );
  
  
  nand q(h, wgaioirl, oezyqhnspy);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [1:1][4:3]  wgaioirl -> logic wgaioirl
  
  not nb(ilvrfefy, oezyqhnspy);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign oezyqhnspy = wgaioirl;
  assign h = 'bx111;
  assign ceegabuwg = '{'{'{'{'bz01,'bz00z0}},'{'{'b10x0x,'bx10x}},'{'{'b1z1,'b0x1}},'{'{'bz0z11,'b01}}},'{'{'{'bzxzx,'bz}},'{'{'b0,'bx}},'{'{'b0xx10,'bxzz}},'{'{'bz01x,'bz}}},'{'{'{'bxzzx,'bz0xxx}},'{'{'bxz1zz,'b1z1x1}},'{'{'b0z,'bz1z}},'{'{'bxz0x,'bz00x}}}};
  assign gbpuekkj = '{'{'bx}};
endmodule: lgogd

module y
  (input bit wyqcmrogg, input trior logic [2:4][3:4][3:0]  ba, input wor logic [4:3] rqysjwzqvk [0:1][0:3][0:1]);
  
  supply1 logic [0:3][2:2][3:4] pkojwqlvp [4:2];
  trireg logic [2:0][4:2][4:4] vpi [2:4][3:0][1:3];
  logic jp [2:4];
  
  xor kbfjhtsk(hhfer, ba, ba);
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   trior logic [2:4][3:4][3:0]  ba -> logic ba
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   trior logic [2:4][3:4][3:0]  ba -> logic ba
  
  not vlc(hhfer, dgy);
  
  lgogd xvvzrhl(.wgaioirl(ba), .ur(jp), .ercrh(vpi), .gbpuekkj(ba), .ceegabuwg(pkojwqlvp));
  // warning: implicit conversion of port connection expands from 2 to 24 bits
  //   logic [1:1][4:3]  wgaioirl -> trior logic [2:4][3:4][3:0]  ba
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   trior logic [2:4][3:4][3:0]  ba -> tri logic [2:2][0:0]  gbpuekkj
  
  not b(ba, dgy);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic ba -> trior logic [2:4][3:4][3:0]  ba
  
  
  // Single-driven assigns
  assign jp = '{'b0x,'b1zzz,'b10zz};
  
  // Multi-driven assigns
  assign ba = wyqcmrogg;
  assign dgy = 'b10000;
endmodule: y

module c
  (output bit aie, output trireg logic [1:3] ldzz [4:0][2:0][2:0], input reg bqdagkrote);
  
  
  
  // Single-driven assigns
  assign aie = aie;
  
  // Multi-driven assigns
endmodule: c

module pmlqvfru
  (output trior logic [2:1][0:0][1:3][4:3] rzpaws [2:2][1:4][4:4][0:3], output wire logic [3:3] hlzfvvzc [1:4][3:4]);
  
  trireg logic [1:3] smebujb [4:0][2:0][2:0];
  
  c bmanzhrypg(.aie(hobqc), .ldzz(smebujb), .bqdagkrote(hnqneho));
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit aie -> wire logic hobqc
  
  nand brnmzn(hnqneho, hnqneho, zh);
  
  not tqvxn(f, jtmgkcsj);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: pmlqvfru



// Seed after: 7659139185679314828,3128299129089410139
