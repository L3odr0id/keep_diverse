// Seed: 9099988925635228673,3128299129089410139

module ljfkte
  (output trireg logic [3:4][0:0][0:4] earc [4:0][3:1][2:4][0:0]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign earc = earc;
endmodule: ljfkte

module duzdyyw
  ( output longint cvnzsno
  , output tri logic [4:0][4:4][0:0] bauageim [3:2]
  , input tri logic [3:4][3:1][2:2] npkbedew [2:0][0:3][3:4][1:4]
  , input tri1 logic palelyr [4:4][3:2][4:0][4:0]
  );
  
  
  
  // Single-driven assigns
  assign cvnzsno = cvnzsno;
  
  // Multi-driven assigns
  assign npkbedew = npkbedew;
  assign palelyr = palelyr;
  assign bauageim = bauageim;
endmodule: duzdyyw

module dgxcdexlvn
  ( output bit [2:3][1:4][1:4][2:0]  g
  , input uwire logic [4:2][2:0][4:4] xsolzxc [4:0]
  , input shortreal hhuoolj
  , input supply1 logic uuvxhzjbd [3:3][0:0][3:3]
  );
  
  trireg logic [3:4][0:0][0:4] rnaub [4:0][3:1][2:4][0:0];
  tri logic [4:0][4:4][0:0] vbwh [3:2];
  tri1 logic hodl [4:4][3:2][4:0][4:0];
  tri logic [3:4][3:1][2:2] gyma [2:0][0:3][3:4][1:4];
  
  duzdyyw xogftoyk(.cvnzsno(g), .bauageim(vbwh), .npkbedew(gyma), .palelyr(hodl));
  // warning: implicit conversion of port connection expands from 64 to 96 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   longint cvnzsno -> bit [2:3][1:4][1:4][2:0]  g
  
  nand nskxsbv(wmdrlyh, g, g);
  // warning: implicit conversion of port connection truncates from 96 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][1:4][1:4][2:0]  g -> logic g
  //
  // warning: implicit conversion of port connection truncates from 96 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][1:4][1:4][2:0]  g -> logic g
  
  ljfkte jwpkbwd(.earc(rnaub));
  
  not hf(wmdrlyh, g);
  // warning: implicit conversion of port connection truncates from 96 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][1:4][1:4][2:0]  g -> logic g
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign gyma = gyma;
  assign wmdrlyh = 'b1;
  assign vbwh = '{'{'{'{'bz}},'{'{'b1zz1z}},'{'{'bxz1x}},'{'{'bz1z}},'{'{'bx}}},'{'{'{'b00x1}},'{'{'b0011}},'{'{'bx11}},'{'{'bz1zz}},'{'{'bz1x10}}}};
  assign hodl = hodl;
endmodule: dgxcdexlvn

module uce
  ( output int rd
  , output tri0 logic [4:3][3:3] vgblnavn [3:3][2:0][2:1]
  , output logic [2:3] lfy [1:1]
  , output triand logic [2:0][4:2][4:3] nhxky [3:3][0:1][1:0][1:4]
  );
  
  
  not kqfik(igpbukmjx, rj);
  
  
  // Single-driven assigns
  assign lfy = lfy;
  assign rd = 'b00;
  
  // Multi-driven assigns
  assign vgblnavn = vgblnavn;
  assign igpbukmjx = rd;
endmodule: uce



// Seed after: 18218363169341951148,3128299129089410139
