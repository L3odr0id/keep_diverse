// Seed: 430576150281111274,3128299129089410139

module ma
  (input bit [2:1][1:3][4:4][2:3]  jf, input reg [2:3] nfowbodnt [3:1][1:2], input bit [3:4]  duj, input bit lto);
  
  
  and yhhy(nl, nl, nl);
  
  not te(nl, nl);
  
  and wqwfalt(nl, duj, lto);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:4]  duj -> logic duj
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit lto -> logic lto
  
  not smlqtfpk(nl, gmp);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign gmp = lto;
endmodule: ma



// Seed after: 18305973876864763085,3128299129089410139
