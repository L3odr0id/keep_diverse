// Seed: 6823947585183604141,3128299129089410139

module c
  (input trireg logic cp [2:1], input integer sc [1:1][1:3], input logic [3:1][1:2]  xjmlpill);
  
  
  nand p(xqafzzmji, xjmlpill, xqafzzmji);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [3:1][1:2]  xjmlpill -> logic xjmlpill
  
  and frbca(lxyionizi, xqafzzmji, lxyionizi);
  
  or iohzv(kgjv, bujmcb, xjmlpill);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [3:1][1:2]  xjmlpill -> logic xjmlpill
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign bujmcb = 'b1;
  assign cp = '{'b0x,'b10};
  assign lxyionizi = xjmlpill;
  assign xqafzzmji = 'b0zz;
endmodule: c

module aaymmqdfn
  (input logic [1:1][0:1][1:3]  eqzixfe, input uwire logic [3:3][2:2][0:3] mxqh [3:2]);
  
  
  nand vwi(ziywwz, uvtxbmcclg, ziywwz);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign uvtxbmcclg = 'b1;
  assign ziywwz = 'b10z;
endmodule: aaymmqdfn

module eqx
  (input trior logic [0:0][3:3]  wognrxbgjy, input trireg logic [2:4][4:0]  agjlfwav);
  
  
  and premcpupaf(fjygacoss, m, m);
  
  and pv(ql, m, m);
  
  not itr(rzr, jxyms);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign m = 'b0zx;
  assign agjlfwav = m;
  assign jxyms = 'b0;
  assign wognrxbgjy = jxyms;
endmodule: eqx



// Seed after: 5245149075574092761,3128299129089410139
