// Seed: 17955976471768091138,3128299129089410139

module xiyda
  ( output real txjxr
  , output bit [1:4][3:1][1:2]  czcd
  , output supply1 logic [2:4] swxwocytu [2:4][0:2][0:1][4:4]
  , output reg [1:4][0:4][4:1] qsj [3:4]
  );
  
  
  nand ffmiuy(czcd, txjxr, t);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic czcd -> bit [1:4][3:1][1:2]  czcd
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real txjxr -> logic txjxr
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign swxwocytu = swxwocytu;
endmodule: xiyda



// Seed after: 11334337321803779299,3128299129089410139
