// Seed: 13510878130923757581,3128299129089410139

module nspoaz
  ( output supply1 logic [3:4] iu [1:2][3:3][1:1]
  , output uwire logic tpxynxpw
  , input supply0 logic [1:1][4:4][1:1] ilox [4:2][0:0][2:4][4:4]
  , input wor logic [2:4][2:2][2:2][2:0] gpjhv [4:3][1:0]
  , input realtime eunnugku
  , input wand logic [1:4][0:2][2:2] zkfspdmme [1:0][3:2]
  );
  
  
  not zlwuyhj(dsvyqbt, gmhuwgcf);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dsvyqbt = tpxynxpw;
  assign gpjhv = gpjhv;
  assign iu = '{'{'{'{'b1x,'bz}}},'{'{'{'bxx0,'bzx0}}}};
  assign zkfspdmme = zkfspdmme;
endmodule: nspoaz

module csgdqb
  ( output tri logic [4:3][1:0] sgwwhw [0:4][2:4][1:3][1:3]
  , output wor logic [2:1][2:2][3:2] jojkjeho [2:0][0:0]
  , output bit [2:4][2:1][0:4]  pve
  , output tri1 logic [1:1] qnb [3:4][0:4][0:4][1:2]
  );
  
  supply1 logic [3:4] uuzypjk [1:2][3:3][1:1];
  wand logic [1:4][0:2][2:2] qdis [1:0][3:2];
  wor logic [2:4][2:2][2:2][2:0] ndoexgf [4:3][1:0];
  supply0 logic [1:1][4:4][1:1] bggdul [4:2][0:0][2:4][4:4];
  
  not qmxvlygpyv(uqi, pve);
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][2:1][0:4]  pve -> logic pve
  
  nand vspp(pve, pve, pve);
  // warning: implicit conversion of port connection expands from 1 to 30 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic pve -> bit [2:4][2:1][0:4]  pve
  //
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][2:1][0:4]  pve -> logic pve
  //
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][2:1][0:4]  pve -> logic pve
  
  nspoaz clqvyfhsf(.iu(uuzypjk), .tpxynxpw(uqi), .ilox(bggdul), .gpjhv(ndoexgf), .eunnugku(pve), .zkfspdmme(qdis));
  // warning: implicit conversion of port connection expands from 30 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][2:1][0:4]  pve -> realtime eunnugku
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign qnb = qnb;
  assign jojkjeho = jojkjeho;
endmodule: csgdqb



// Seed after: 2167559344450510339,3128299129089410139
