// Seed: 5893021453546226726,3128299129089410139

module ugiqt
  (input trireg logic [2:4][4:1]  kyu, input supply1 logic [1:4][4:2] igyb [3:1][3:2][1:2]);
  
  
  and ysu(kyu, kyu, kyu);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic kyu -> trireg logic [2:4][4:1]  kyu
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   trireg logic [2:4][4:1]  kyu -> logic kyu
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   trireg logic [2:4][4:1]  kyu -> logic kyu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ugiqt



// Seed after: 5099076482301640435,3128299129089410139
