// Seed: 8966281038822525192,3128299129089410139

module naplhcsfn
  ( output byte bqpqf
  , output time c
  , output reg raczpwte [1:0][2:2]
  , input wand logic [1:2][2:4][2:2] qevqinxh [3:0]
  , input uwire logic aadmvw [3:4][1:4][0:4][3:0]
  );
  
  
  nand uw(wyupflmo, wyupflmo, kt);
  
  
  // Single-driven assigns
  assign bqpqf = wyupflmo;
  assign c = bqpqf;
  
  // Multi-driven assigns
endmodule: naplhcsfn



// Seed after: 6580800625636262848,3128299129089410139
