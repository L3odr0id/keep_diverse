// Seed: 3253010377385789457,3128299129089410139

module wwpfdexi
  (output logic [4:2][1:0][2:2][0:2]  tragboep, output int dxsakpnwc);
  
  
  
  // Single-driven assigns
  assign tragboep = '{'{'{'{'bx0,'bzzx,'b1xx01}},'{'{'b0,'bz11,'b1xz}}},'{'{'{'bx0zz,'b0xz0,'b1xxx}},'{'{'bxz111,'bz1,'bx}}},'{'{'{'b1x,'b01,'bz}},'{'{'bz01z0,'bzz0xx,'bz1}}}};
  assign dxsakpnwc = 'b1101;
  
  // Multi-driven assigns
endmodule: wwpfdexi



// Seed after: 12506491258351115114,3128299129089410139
