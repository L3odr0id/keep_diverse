// Seed: 15066836924594815433,3128299129089410139

module ltfgm
  ( output reg [1:3]  wdinqy
  , output reg [0:2]  pblaxm
  , output reg [0:1][0:2][4:1]  iwskafltk
  , output supply1 logic [1:0][0:0][2:1]  bkpagblwf
  , input trior logic [1:1] i [0:2][3:3][0:3][1:2]
  , input trireg logic [4:1] lbxjjsjbzm [1:2][1:1][1:4][3:1]
  );
  
  
  
  // Single-driven assigns
  assign wdinqy = '{'bz0xxx,'b0,'b1zx1};
  assign iwskafltk = '{'{'{'b1xx0,'b1xz,'b1z00x,'b1},'{'bz0110,'b0,'b011,'b11x},'{'b1xx1,'b10,'bxx11,'b0}},'{'{'bx,'b0z11,'bz,'bzxxx0},'{'bx0xz,'bxz110,'b0010x,'bzzzx},'{'bzz,'bz,'b10zx,'bxzzz1}}};
  assign pblaxm = iwskafltk;
  
  // Multi-driven assigns
endmodule: ltfgm

module f
  ( output bit uuihh
  , input trior logic [3:3][1:2] ffwya [3:4]
  , input shortreal fbelcrnkh
  , input trireg logic [3:1] enoj [4:3][3:0][0:1]
  , input supply1 logic j [1:3][4:4][2:3]
  );
  
  
  or semhrwsp(uuihh, uuihh, fbelcrnkh);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic uuihh -> bit uuihh
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit uuihh -> logic uuihh
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal fbelcrnkh -> logic fbelcrnkh
  
  not rpqvumtco(vsqt, fbelcrnkh);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal fbelcrnkh -> logic fbelcrnkh
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ffwya = ffwya;
  assign enoj = enoj;
endmodule: f

module ambnl
  ( output tri logic q [3:1][4:1][0:3]
  , output reg [0:2]  nnwpianaqi
  , output logic a [0:0]
  , input logic d
  , input logic [3:2][0:1][3:0] oyleueq [4:4]
  );
  
  
  
  // Single-driven assigns
  assign nnwpianaqi = '{'bzx,'bx,'bzz0xz};
  assign a = a;
  
  // Multi-driven assigns
  assign q = q;
endmodule: ambnl

module k
  ( output logic [3:3][3:1][3:1][1:3]  tvsbswur
  , output triand logic [4:4][4:4]  hgixjjnnn
  , input longint yuvoofcviu
  , input bit [1:3][2:0] xilbsnhld [2:0][2:1]
  , input bit n
  );
  
  
  
  // Single-driven assigns
  assign tvsbswur = '{'{'{'{'b0z1,'bzz,'bxxx},'{'bxx1xx,'b1x1zz,'bx},'{'bxxx0,'b11x,'b10x}},'{'{'b0zzx1,'bx0z1,'bx0},'{'b0z111,'bzx,'b10z},'{'bx0x,'bz1,'b011x}},'{'{'b1x00x,'b1,'b11},'{'b1x0x,'bxx1,'bz},'{'b0zz,'bz000,'b100}}}};
  
  // Multi-driven assigns
  assign hgixjjnnn = '{'{'b1z11}};
endmodule: k



// Seed after: 16755045049282625894,3128299129089410139
