// Seed: 11800529220501756588,3128299129089410139

module vetujnovpx
  ( output bit [1:3][3:1][4:0]  khmrgsehz
  , input int jchpzv
  , input supply0 logic [0:0] gebnt [4:4][4:3][4:1][1:0]
  , input supply0 logic [4:4][3:1]  sw
  );
  
  
  and vxd(khmrgsehz, re, lmkvo);
  // warning: implicit conversion of port connection expands from 1 to 45 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic khmrgsehz -> bit [1:3][3:1][4:0]  khmrgsehz
  
  and jipxwucp(lmkvo, ukmgjepdgf, re);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign re = 'b1;
  assign gebnt = gebnt;
  assign ukmgjepdgf = 'b0;
  assign lmkvo = lmkvo;
endmodule: vetujnovpx

module fssq
  (output logic fmb [0:0], output logic [4:3] lgwtsl [1:1][0:2], output wand logic [3:3][4:0] qhtrsnvven [2:2][1:1]);
  
  
  
  // Single-driven assigns
  assign lgwtsl = '{'{'{'b01,'bx00z},'{'bz1x1z,'b1x1},'{'bxzx0x,'b10z}}};
  assign fmb = '{'bz1};
  
  // Multi-driven assigns
  assign qhtrsnvven = '{'{'{'{'bzz,'b11,'b00xxx,'b0,'b00}}}};
endmodule: fssq



// Seed after: 2519640146387862472,3128299129089410139
