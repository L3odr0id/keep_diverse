// Seed: 9407371298728588963,3128299129089410139

module bcn
  (output supply1 logic [2:1][0:1] fuox [2:3][4:4][0:3]);
  
  
  not lseaqk(kdtgkge, kdtgkge);
  
  or xqnxukq(kdtgkge, cwi, y);
  
  or dgcffyy(leexct, cwi, bmcd);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kdtgkge = leexct;
  assign bmcd = kdtgkge;
  assign y = 'b0x1z;
  assign cwi = bmcd;
  assign fuox = fuox;
endmodule: bcn



// Seed after: 7958188861447328083,3128299129089410139
