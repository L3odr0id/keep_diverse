// Seed: 18218363169341951148,3128299129089410139

module cvjqrwm
  ( output uwire logic [1:3][3:2] jq [3:2][0:2][0:2]
  , output reg szrxjwmj
  , output shortint ivi [1:2]
  , output tri logic [1:4][2:0][4:1][3:4]  fqyxdnf
  , input reg [2:0][1:1][2:0][0:2]  jfe
  , input reg [1:4]  ygl
  , input logic [4:0]  xcxn
  );
  
  
  not yexelc(hcokdbtjgg, szrxjwmj);
  
  
  // Single-driven assigns
  assign szrxjwmj = jfe;
  assign jq = jq;
  
  // Multi-driven assigns
  assign fqyxdnf = '{'{'{'{'b0x1,'b0},'{'bx00,'bx01},'{'b0x,'bz101},'{'bz101,'b1x}},'{'{'b1,'b10z},'{'b01zx,'bx10},'{'b01,'bx00},'{'bz0z1,'b1zz}},'{'{'b11x,'b11xx},'{'bz1xz,'b11zzz},'{'b0x01z,'bx11z0},'{'bx0zx1,'bz}}},'{'{'{'bx11x,'b111x},'{'b11x,'b1x10z},'{'b0x0x0,'b0},'{'b1010z,'bx01x0}},'{'{'bz,'bz01},'{'bz00x,'b0100},'{'bz,'b0},'{'bxz0xz,'bxz}},'{'{'bxx1xx,'b1},'{'bz0,'b1z11},'{'b1z,'bzx},'{'b0,'bz01x1}}},'{'{'{'b1101,'bx1},'{'b1x00z,'bxx},'{'bxx0,'b0zxz},'{'b00xxx,'b0x}},'{'{'b010z,'bz100},'{'b111,'b01},'{'b0,'b11x0},'{'b1xxx,'b1x0zz}},'{'{'bx110x,'b010xx},'{'bx10z,'b00x},'{'bz01,'b11},'{'bz11,'bz11}}},'{'{'{'bx00,'bx0001},'{'b00z,'bx0xx},'{'b00z0z,'b0xx},'{'b1x111,'b01x}},'{'{'bz,'bz},'{'bxz,'b0x0z1},'{'b1,'b1xzx0},'{'b1,'bzz0z}},'{'{'bz,'b001},'{'bx,'bz1},'{'b10x,'bzxx10},'{'bxx,'b1010}}}};
  assign hcokdbtjgg = 'bz;
endmodule: cvjqrwm

module cmmo
  (input reg [0:1][0:3][1:0]  y, input logic [4:2][4:3]  sra);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: cmmo

module cysiq
  ( input trireg logic [2:0][4:1] dmpqgs [0:4][2:4][1:3][3:4]
  , input trireg logic [3:1][1:3][2:0][3:4] rlzksilyyo [2:4][2:0][3:1]
  , input logic [2:3][4:4][4:3][3:2]  anot
  );
  
  
  nand wgcfqronad(hfw, luimluusjy, luimluusjy);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rlzksilyyo = rlzksilyyo;
  assign dmpqgs = dmpqgs;
  assign luimluusjy = 'bx;
endmodule: cysiq



// Seed after: 3117070915413338426,3128299129089410139
