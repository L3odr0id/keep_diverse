// Seed: 3117070915413338426,3128299129089410139

module m
  ( output wire logic [2:4][3:2]  rrwzikdx
  , output reg [0:3][4:0]  jop
  , output wire logic [3:2] w [4:3][0:2]
  , output reg [4:1] evzkzb [0:3]
  , input bit mhhpm [2:2]
  );
  
  
  or xudi(gxow, rrwzikdx, rrwzikdx);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   wire logic [2:4][3:2]  rrwzikdx -> logic rrwzikdx
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   wire logic [2:4][3:2]  rrwzikdx -> logic rrwzikdx
  
  xor obzi(cs, rrwzikdx, jop);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   wire logic [2:4][3:2]  rrwzikdx -> logic rrwzikdx
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   reg [0:3][4:0]  jop -> logic jop
  
  and birzuhqh(e, cs, okdn);
  
  not arsv(kgll, ioehh);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ioehh = gxow;
  assign gxow = 'b1z0z;
  assign w = '{'{'{'b0,'bz00},'{'b11z,'bzx0zz},'{'bx0,'b1}},'{'{'bx0,'b1},'{'b1,'b1x11x},'{'bzx,'bz100z}}};
  assign rrwzikdx = rrwzikdx;
endmodule: m

module rz
  (output logic [2:0][4:1][3:1]  tpw, output uwire logic [0:3][1:3] obybcea [4:3][4:2][4:1][3:1]);
  
  
  or whvsb(b, tpw, tpw);
  // warning: implicit conversion of port connection truncates from 36 to 1 bits
  //   logic [2:0][4:1][3:1]  tpw -> logic tpw
  //
  // warning: implicit conversion of port connection truncates from 36 to 1 bits
  //   logic [2:0][4:1][3:1]  tpw -> logic tpw
  
  not ely(tpw, r);
  // warning: implicit conversion of port connection expands from 1 to 36 bits
  //   logic tpw -> logic [2:0][4:1][3:1]  tpw
  
  
  // Single-driven assigns
  assign obybcea = obybcea;
  
  // Multi-driven assigns
endmodule: rz

module xkmmrmcufl
  (output int thxjrx [4:2], input bit [1:1][3:1] w [3:0]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: xkmmrmcufl



// Seed after: 11532771568697646238,3128299129089410139
