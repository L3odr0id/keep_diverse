// Seed: 15337481340297115087,3128299129089410139

module folvob
  (output reg [2:2][4:3][4:3][0:2]  oqkfdauat, input trireg logic [3:4][1:3][0:1][0:2]  jp);
  
  
  nand cmc(oqkfdauat, ngpppre, wjr);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic oqkfdauat -> reg [2:2][4:3][4:3][0:2]  oqkfdauat
  
  or jxy(jp, wvabgkxsn, rtafefzawk);
  // warning: implicit conversion of port connection expands from 1 to 36 bits
  //   logic jp -> trireg logic [3:4][1:3][0:1][0:2]  jp
  
  not dbuwvmmezx(z, zqbswmoeec);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ngpppre = oqkfdauat;
  assign jp = '{'{'{'{'bx1,'bz,'bz},'{'b1,'bx,'bzz}},'{'{'bxz00,'b1zx,'bz},'{'bz0,'bx0,'bx}},'{'{'b1,'bxz01,'b01},'{'bx0,'bx1,'b0}}},'{'{'{'b0zz,'bxzzxx,'b11},'{'bxx0z,'b11,'b1z11}},'{'{'bzx0zx,'b0001z,'b1x},'{'b1x1z,'bzxx0,'b0}},'{'{'bx10zx,'bxxxx,'b0x},'{'b10x01,'bx,'bz1}}}};
  assign wvabgkxsn = 'bz;
  assign rtafefzawk = 'bzxxx1;
  assign wjr = wjr;
endmodule: folvob

module x
  ( output bit [1:4][1:0]  s
  , output reg [1:0] jbpimbc [2:3]
  , output bit pvw
  , output bit [3:2][2:4]  q
  , input tri1 logic [1:1] sc [0:3][1:2][3:4]
  , input trireg logic [4:1][2:4]  sqazqrclv
  );
  
  
  
  // Single-driven assigns
  assign s = '{'{'b1111,'b0000},'{'b0,'b11},'{'b101,'b0111},'{'b0,'b00100}};
  
  // Multi-driven assigns
  assign sqazqrclv = '{'{'b11x1x,'bx,'bz00z},'{'bx,'bx10,'bx},'{'bz1xz1,'bxz,'bx1x0x},'{'bzx,'b01x,'b01x}};
endmodule: x

module fq
  (output bit sypqine [1:1], input wire logic [2:1][3:0]  wxodyq, input uwire logic [4:4] ieanca [3:1][2:4]);
  
  
  
  // Single-driven assigns
  assign sypqine = sypqine;
  
  // Multi-driven assigns
  assign wxodyq = wxodyq;
endmodule: fq



// Seed after: 17120606345259600647,3128299129089410139
