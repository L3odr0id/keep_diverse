// Seed: 13647994075863507267,3128299129089410139

module vsmopgmv
  ( output bit [2:0][1:2][1:3]  poy
  , output longint vhcfoqerv [1:0][4:3]
  , output bit [0:0][0:3][2:4] pvkgowgx [3:0]
  , input tri0 logic [2:3][4:2][3:4][0:3] nlpqdkywom [2:4][0:1]
  , input tri logic [0:0][2:0][0:2] s [2:2]
  );
  
  
  not cz(poy, poy);
  // warning: implicit conversion of port connection expands from 1 to 18 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic poy -> bit [2:0][1:2][1:3]  poy
  //
  // warning: implicit conversion of port connection truncates from 18 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:0][1:2][1:3]  poy -> logic poy
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nlpqdkywom = nlpqdkywom;
  assign s = s;
endmodule: vsmopgmv



// Seed after: 328071024425920796,3128299129089410139
