// Seed: 12475482197253238135,3128299129089410139

module ocebcv
  ( output supply0 logic [2:0] ylx [1:0][4:4][0:2]
  , output wor logic [4:1][3:4][4:2][1:2] evwtpbzg [0:4][2:3]
  , input reg [1:3] swxcgzpwa [1:4]
  , input reg lamxtds [1:2]
  , input reg [2:4][3:0]  kctkr
  , input uwire logic ljrrjmunf [2:3]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ylx = ylx;
  assign evwtpbzg = evwtpbzg;
endmodule: ocebcv



// Seed after: 3253010377385789457,3128299129089410139
