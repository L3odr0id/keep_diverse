// Seed: 4730330285713594232,3128299129089410139

module uqcckhdj
  ( output reg [0:2][3:3]  kzrbtozob
  , input wor logic [3:2][3:1]  fm
  , input triand logic pjl [3:0][3:0][1:0]
  , input reg [1:2][0:2] xsjyrdc [2:1][4:2]
  , input int sw
  );
  
  
  xor qxwxaiqtc(kzrbtozob, kzrbtozob, kzrbtozob);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic kzrbtozob -> reg [0:2][3:3]  kzrbtozob
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][3:3]  kzrbtozob -> logic kzrbtozob
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][3:3]  kzrbtozob -> logic kzrbtozob
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: uqcckhdj



// Seed after: 5555284318056057502,3128299129089410139
