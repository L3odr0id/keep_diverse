// Seed: 15791412969388589653,3128299129089410139

module yvjdma
  ( output supply0 logic [2:2][0:2][1:4][0:1] ulbq [3:4][4:4][3:4]
  , output wire logic [0:4]  wvk
  , input supply1 logic [4:4][1:1][0:4] l [2:0][4:3]
  , input logic [4:0][2:1]  xhcwlcju
  );
  
  
  nand dclvaxgnkf(mspsjr, cwczfkhv, odrkf);
  
  xor fisquafey(foiexehwih, wvk, cwczfkhv);
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   wire logic [0:4]  wvk -> logic wvk
  
  not v(oayb, jojoa);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign l = l;
  assign wvk = foiexehwih;
  assign ulbq = ulbq;
  assign jojoa = 'bz;
  assign oayb = wvk;
endmodule: yvjdma

module o
  (input logic [3:0] bawwr [1:1][1:1], input bit twl [0:3], input wand logic ethmvhrrft, input trireg logic [1:0][3:2] alrfg [0:3]);
  
  
  and cwdhoik(ulgq, ethmvhrrft, bvslsx);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ethmvhrrft = 'b0zz0x;
  assign bvslsx = ethmvhrrft;
endmodule: o



// Seed after: 1148233422042294380,3128299129089410139
