// Seed: 4261191817767376468,3128299129089410139

module lzfrlvv
  (input tri0 logic [4:2][3:4][3:1][3:1]  rliyyh, input realtime iwayhse, input reg [3:0] fnkbbd [0:4]);
  
  
  not fefxrqihgk(nffsjkhwj, dp);
  
  not ppchjzizr(gjnjdgurf, virzhti);
  
  not ldajhlrrj(s, lexf);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign s = 'b1x;
  assign virzhti = iwayhse;
  assign rliyyh = '{'{'{'{'b10z00,'b0zxx0,'b1},'{'b00,'bzzx,'bxzxzz},'{'bzxxx,'bz,'b00xzx}},'{'{'bz0,'b1zx,'b0x1},'{'bzz00,'b001z,'bzxz1z},'{'bz10z,'bx,'bz1zx1}}},'{'{'{'b10,'b0xx,'b1},'{'b0x,'bz01,'bx1},'{'b0x11,'b001x,'bzz}},'{'{'bxxxx,'b0,'b0},'{'bxx1,'b1,'b0x},'{'b1zz0,'bx11xx,'b10x1x}}},'{'{'{'bxz1x,'bz110,'b10z},'{'b0zx,'b1xxz,'bz},'{'bxz,'b0,'bzx0z}},'{'{'bx00x0,'bx,'b0xz},'{'b0zzx,'b010,'b1xz},'{'bxz,'bzx0,'bzz1z1}}}};
  assign dp = 'b010x;
  assign lexf = dp;
endmodule: lzfrlvv

module ktaryq
  ( input supply0 logic [1:3][3:0]  jz
  , input reg [0:0][2:0]  oja
  , input supply1 logic wh [3:1][3:4]
  , input supply0 logic [2:4][0:3][0:2] creo [1:0][2:4]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign creo = creo;
  assign wh = '{'{'bx11zz,'bx100z},'{'b0,'b111},'{'b0z11x,'b0}};
  assign jz = '{'{'bx110x,'bz011z,'bz,'b111},'{'b11100,'bzx1z1,'b11z1,'bz1},'{'bzxzz0,'b1x0z,'bxz1z,'b1x1}};
endmodule: ktaryq



// Seed after: 7075531678909538591,3128299129089410139
