// Seed: 5099076482301640435,3128299129089410139

module fweczzumxf
  ( input uwire logic [1:1][1:0] htentqieap [0:0]
  , input uwire logic [2:0][3:4] uguu [4:0][0:1][1:0]
  , input bit [3:1][0:2][1:3][4:3]  fycry
  , input reg [0:4][3:2]  hnvfopc
  );
  
  
  not ehridfpwbb(rz, jp);
  
  xor rmydfuk(rpguagdaab, nwsc, svpkwmvkzb);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rpguagdaab = rpguagdaab;
  assign jp = 'bx0z11;
  assign nwsc = nwsc;
endmodule: fweczzumxf

module bzmowyad
  (output byte kdboh [4:0][4:1], output longint ggbeyfhuz, output wire logic [1:2][3:4]  qbscc);
  
  
  not xyoirnx(ggbeyfhuz, ggbeyfhuz);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic ggbeyfhuz -> longint ggbeyfhuz
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ggbeyfhuz -> logic ggbeyfhuz
  
  nand rwvubplcml(bbzjwpxde, mh, bbzjwpxde);
  
  not zhnmpeeeoh(bqohwjyw, lypmeffgg);
  
  xor ecxvwgwqar(ubl, bbzjwpxde, lypmeffgg);
  
  
  // Single-driven assigns
  assign kdboh = kdboh;
  
  // Multi-driven assigns
  assign mh = ubl;
endmodule: bzmowyad

module jcqvzdtis
  ( output reg atrgzhzf
  , output bit [3:3] nks [1:3][1:3]
  , output wire logic [0:4][2:1][0:4][3:1] fnd [1:0][1:2]
  , input uwire logic [1:2][2:0][2:2][4:2] vxfyico [0:2]
  , input tri logic [1:2][0:0] qso [4:1]
  , input longint rgjd
  , input trior logic [3:2] hrx [0:4][0:4][4:2][2:4]
  );
  
  
  not zp(atrgzhzf, rgjd);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint rgjd -> logic rgjd
  
  xor f(qofb, assqwow, assqwow);
  
  
  // Single-driven assigns
  assign nks = nks;
  
  // Multi-driven assigns
endmodule: jcqvzdtis



// Seed after: 13647994075863507267,3128299129089410139
