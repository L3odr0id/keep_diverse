// Seed: 12658144569597683733,3128299129089410139

module imlsl
  ( output wor logic [2:4][1:1]  k
  , output bit igrwyabbjl [4:4][4:4]
  , output trireg logic [4:3]  xosnvbkr
  , output reg [0:3][2:1][1:4]  evsucutd
  , input wor logic [4:2][4:2] eeg [4:1][4:3][3:2][3:0]
  , input shortreal vr
  , input triand logic [1:4][0:2] kbfxv [2:1][3:0][0:2][3:4]
  , input bit [1:1][3:0][2:4] xxdcf [2:3]
  );
  
  
  and oiwx(aplesvy, vr, k);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal vr -> logic vr
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wor logic [2:4][1:1]  k -> logic k
  
  not tnwtjqesc(xgfpgtsj, nyfgllfayh);
  
  not hwutqobmpy(xtqobpoc, rplvxnqej);
  
  
  // Single-driven assigns
  assign igrwyabbjl = '{'{'b0010}};
  assign evsucutd = k;
  
  // Multi-driven assigns
  assign xosnvbkr = xosnvbkr;
  assign nyfgllfayh = 'bxzxz0;
  assign rplvxnqej = k;
endmodule: imlsl

module orfhsx
  (output reg pbnvqcc, output wor logic [1:3][4:3][2:0][3:3] fw [3:0][4:0][0:2][4:2], output reg u, input shortint rth);
  
  bit pg [4:4][4:4];
  bit [1:1][3:0][2:4] ului [2:3];
  triand logic [1:4][0:2] iylhzxmq [2:1][3:0][0:2][3:4];
  wor logic [4:2][4:2] hrlv [4:1][4:3][3:2][3:0];
  
  nand lvhmip(qrcd, tq, pbnvqcc);
  
  nand y(u, dyyibwrdg, pbnvqcc);
  
  imlsl fvandlf(.k(rdlakooqha), .igrwyabbjl(pg), .xosnvbkr(ewfytglvx), .evsucutd(s), .eeg(hrlv), .vr(hlj), .kbfxv(iylhzxmq), .xxdcf(ului));
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wor logic [2:4][1:1]  k -> wire logic rdlakooqha
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   trireg logic [4:3]  xosnvbkr -> wire logic ewfytglvx
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   reg [0:3][2:1][1:4]  evsucutd -> wire logic s
  //
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic hlj -> shortreal vr
  
  or yurgoayzrc(pbnvqcc, rth, u);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint rth -> logic rth
  
  
  // Single-driven assigns
  assign ului = '{'{'{'{'b010,'b01001,'b101},'{'b111,'b0110,'b001},'{'b00,'b0,'b11},'{'b0,'b1001,'b000}}},'{'{'{'b1100,'b0100,'b0},'{'b10,'b1011,'b00100},'{'b1101,'b011,'b01100},'{'b11,'b10,'b1}}}};
  
  // Multi-driven assigns
  assign rdlakooqha = ewfytglvx;
  assign dyyibwrdg = dyyibwrdg;
  assign fw = fw;
endmodule: orfhsx

module yzswrw
  (output tri logic [0:0] oeihwitsab [3:1][4:4][0:1][3:1]);
  
  
  or drdl(yyzercxr, yyzercxr, wlmckp);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign oeihwitsab = oeihwitsab;
  assign yyzercxr = wlmckp;
  assign wlmckp = 'b011zz;
endmodule: yzswrw

module whunoj
  ( input trior logic [0:1][2:2][4:4][2:3] olnw [3:1][0:0]
  , input triand logic lfstqjbmfi [2:1][4:4][1:3][3:2]
  , input bit [0:4][2:3]  ql
  , input wor logic [2:4][1:1][2:4][2:2] trhyhczc [4:3][0:1][1:3]
  );
  
  wor logic [1:3][4:3][2:0][3:3] lrtbxmepo [3:0][4:0][0:2][4:2];
  
  nand ezcjgvj(xnymgk, xnymgk, yo);
  
  and vng(xnymgk, vrlljmvhw, xnymgk);
  
  and zmci(npggrzqnx, mf, yo);
  
  orfhsx dhzh(.pbnvqcc(oks), .fw(lrtbxmepo), .u(cqhpb), .rth(vrlljmvhw));
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic vrlljmvhw -> shortint rth
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xnymgk = 'b11;
  assign vrlljmvhw = 'bzzz1x;
  assign npggrzqnx = 'bx;
  assign yo = xnymgk;
endmodule: whunoj



// Seed after: 10303539322999713515,3128299129089410139
