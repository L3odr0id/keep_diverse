// Seed: 4773139017576541913,3128299129089410139

module camchgxb
  ( output tri logic [0:3] dxsfriimm [1:3][3:3]
  , output bit wudixi [0:4]
  , output triand logic [2:3][0:1] lvrgtkp [3:3][4:4][4:4][1:2]
  , input supply1 logic hd [0:4]
  , input wire logic [4:0] isdkd [1:2][4:0]
  , input tri1 logic [4:3] rbxvpoo [2:1][0:0]
  , input bit [4:3][2:4]  t
  );
  
  
  nand gt(ulai, ulai, ulai);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rbxvpoo = rbxvpoo;
  assign lvrgtkp = lvrgtkp;
  assign dxsfriimm = dxsfriimm;
endmodule: camchgxb

module qylvl
  ( output wire logic [0:4][0:0][0:2] nszhsash [3:4][1:4][3:1]
  , input logic zyu
  , input trior logic [2:4][3:3][1:3] hwej [1:0]
  , input triand logic [0:2]  viirnxmvcj
  );
  
  
  xor fxtli(viirnxmvcj, zyu, zyu);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic viirnxmvcj -> triand logic [0:2]  viirnxmvcj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nszhsash = nszhsash;
  assign hwej = '{'{'{'{'b0z0z,'b1,'bx00}},'{'{'b1xx1,'b0,'b1z1x}},'{'{'b01,'bx,'b01}}},'{'{'{'bxz0zz,'b0z,'b0x}},'{'{'b000,'bz1zz0,'bxzzx}},'{'{'b00,'b1zxz1,'bz1x}}}};
endmodule: qylvl



// Seed after: 15066836924594815433,3128299129089410139
