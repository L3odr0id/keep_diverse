// Seed: 13299826562397828311,3128299129089410139

module fc
  (output supply1 logic [1:0][4:1][0:2][4:4] mrucan [4:1][4:3][0:2], input tri0 logic [2:0][0:0][1:2] gxhyhkraf [4:2], input bit tce);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign mrucan = mrucan;
  assign gxhyhkraf = gxhyhkraf;
endmodule: fc

module ye
  ( output supply0 logic [2:3] jwqf [1:1][2:3]
  , output trireg logic rbpljgp [4:1]
  , input supply0 logic [1:1][4:2][4:0] r [1:4][4:1][0:0][1:2]
  , input triand logic [0:1][1:4][0:0][0:4] tjmgok [2:3][1:1][3:3]
  );
  
  supply1 logic [1:0][4:1][0:2][4:4] suxb [4:1][4:3][0:2];
  tri0 logic [2:0][0:0][1:2] laenbfcf [4:2];
  
  nand fzrtwe(a, arkuy, hzffa);
  
  fc n(.mrucan(suxb), .gxhyhkraf(laenbfcf), .tce(t));
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic t -> bit tce
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign a = arkuy;
  assign hzffa = t;
endmodule: ye

module qyipbxecf
  ( output reg jcdg
  , output reg g
  , output triand logic [4:3][1:3] pknbi [0:0][3:2]
  , input reg [0:3] eskjwd [2:0]
  , input tri1 logic [1:1]  uupemuncj
  , input triand logic bce [4:4]
  , input trior logic [0:0][3:0][2:0] xxllkir [0:2]
  );
  
  
  or mkehuri(b, bvhxhjabu, bmbr);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign b = jcdg;
  assign uupemuncj = jcdg;
  assign bvhxhjabu = 'b0zxx;
  assign bmbr = jcdg;
endmodule: qyipbxecf

module igbxcw
  ( output tri1 logic [3:0] tnynbqge [1:3][1:1][4:3][0:4]
  , output trireg logic [0:0][1:4][2:2][0:0] hrkfnh [4:0][0:1]
  , input wor logic [1:2][2:1] ufw [1:2][4:2][4:1]
  , input triand logic [3:3][3:1][0:3] xyj [3:3][3:4][1:1]
  , input reg [0:3]  qg
  );
  
  
  xor lfgrp(alszltw, jv, jwbml);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: igbxcw



// Seed after: 2775971243336691657,3128299129089410139
