// Seed: 8355443864916960300,3128299129089410139

module euol
  (output logic [4:1][1:3][1:4][2:3]  x, output reg [1:2][3:4][3:0]  hoe);
  
  
  not ihxzpt(x, hoe);
  // warning: implicit conversion of port connection expands from 1 to 96 bits
  //   logic x -> logic [4:1][1:3][1:4][2:3]  x
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   reg [1:2][3:4][3:0]  hoe -> logic hoe
  
  or yyr(hoe, hoe, x);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  //   logic hoe -> reg [1:2][3:4][3:0]  hoe
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   reg [1:2][3:4][3:0]  hoe -> logic hoe
  //
  // warning: implicit conversion of port connection truncates from 96 to 1 bits
  //   logic [4:1][1:3][1:4][2:3]  x -> logic x
  
  or sunb(iutlan, hoe, w);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   reg [1:2][3:4][3:0]  hoe -> logic hoe
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: euol

module hpdnjj
  ( output supply0 logic uhptkf
  , output real wavyccrs
  , input logic [2:1][2:0][0:3][1:2]  y
  , input wire logic [3:3] hpyddad [2:4]
  , input trior logic [0:2][0:0][3:0] qhnsu [4:2]
  );
  
  
  or xmo(pxouvqoham, uhptkf, uhptkf);
  
  
  // Single-driven assigns
  assign wavyccrs = y;
  
  // Multi-driven assigns
  assign qhnsu = '{'{'{'{'bz0,'b11x00,'b01x,'b0}},'{'{'b00z01,'b1,'bxzx1z,'bz00z}},'{'{'bx0,'bx001,'b1z10,'b0xz}}},'{'{'{'bz,'bz,'b1z10,'b0}},'{'{'bzz0,'bx,'b00x01,'bxx}},'{'{'bxzx,'bz01,'bz0,'b10xx}}},'{'{'{'bxz0,'b11z0,'bxz,'bxxx1}},'{'{'b0xzx,'b1,'b1001,'b1}},'{'{'b0,'b0,'b0x,'b000x}}}};
  assign uhptkf = uhptkf;
  assign pxouvqoham = 'b1z1;
endmodule: hpdnjj

module eusn
  (output trior logic [3:3][1:3] saxtswwhk [2:0], output reg kbu, input triand logic [1:4] sxodqqfbzf [1:1][1:1], input logic lnkgzte);
  
  
  euol rgrakx(.x(kbu), .hoe(dvdxpndqj));
  // warning: implicit conversion of port connection truncates from 96 to 1 bits
  //   logic [4:1][1:3][1:4][2:3]  x -> reg kbu
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   reg [1:2][3:4][3:0]  hoe -> wire logic dvdxpndqj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign sxodqqfbzf = sxodqqfbzf;
endmodule: eusn



// Seed after: 1536635323995096370,3128299129089410139
