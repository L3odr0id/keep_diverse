// Seed: 1735739043436887574,3128299129089410139

module qlg
  (input wand logic [3:3] ihhcjw [0:4][4:3], input bit kew, input bit [2:1][4:3][3:3][3:3]  wmilyybbn, input real rlwcseg [2:3]);
  
  
  not hy(gol, vyxfx);
  
  not lurj(vyxfx, vyxfx);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign vyxfx = 'bzz1;
  assign ihhcjw = '{'{'{'bx1z0x},'{'bx1}},'{'{'b110z},'{'b01z}},'{'{'b1z01z},'{'b1xz}},'{'{'bx0x},'{'bz10z1}},'{'{'bx},'{'bx0z0}}};
endmodule: qlg



// Seed after: 10452617400833083778,3128299129089410139
