// Seed: 13966551278677208945,3128299129089410139

module xgvwfo
  ( output wor logic [3:3][0:3]  xwvmwksxo
  , output tri1 logic aqq [4:1][3:1][4:2]
  , input trireg logic [0:2] piemvgww [1:0][1:2]
  , input bit [0:1][2:4][0:2] asseuoeqd [3:0]
  , input wor logic [0:0] jruhfmtat [1:3][2:0]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: xgvwfo

module iiprng
  ( output triand logic [2:2][4:2][3:4] ggvggpjabh [1:3][4:4][0:0]
  , output logic ckc [0:4]
  , output supply0 logic [4:2][4:3] lml [2:2]
  , input logic [1:3][3:2][0:3]  gtrzosmn
  );
  
  
  or lbc(egw, gtrzosmn, gtrzosmn);
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   logic [1:3][3:2][0:3]  gtrzosmn -> logic gtrzosmn
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   logic [1:3][3:2][0:3]  gtrzosmn -> logic gtrzosmn
  
  
  // Single-driven assigns
  assign ckc = ckc;
  
  // Multi-driven assigns
  assign egw = 'b0x1;
  assign lml = lml;
  assign ggvggpjabh = ggvggpjabh;
endmodule: iiprng



// Seed after: 17571190611611453888,3128299129089410139
