// Seed: 7659139185679314828,3128299129089410139

module ntfsx
  ( output reg [0:4][3:1][3:3] lslarkfyv [0:2]
  , output trior logic [0:4][3:0][4:1][0:2] muyhuoih [1:0][3:0][4:0][1:3]
  , output shortreal t
  , output realtime btb
  , input realtime kv
  , input tri1 logic [0:0][1:4][0:4][0:2] ticxteghen [3:3]
  , input tri logic [0:3][1:1][3:4][1:0] vlfuhut [3:3]
  , input wand logic [2:4][4:0]  bss
  );
  
  
  nand a(t, t, t);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic t -> shortreal t
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal t -> logic t
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal t -> logic t
  
  and d(drqqy, btb, huqww);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime btb -> logic btb
  
  not njdc(nrvup, t);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal t -> logic t
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign drqqy = 'b00x;
  assign ticxteghen = ticxteghen;
  assign nrvup = 'b000z0;
  assign vlfuhut = vlfuhut;
  assign muyhuoih = muyhuoih;
endmodule: ntfsx

module wvmtb
  (output bit mrcyxwzl [0:3][1:1][2:2], output longint eovcuyo, output reg [4:3] lns [3:1]);
  
  
  not uuj(eovcuyo, eovcuyo);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic eovcuyo -> longint eovcuyo
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint eovcuyo -> logic eovcuyo
  
  xor wir(syferkh, hbfehdouq, syferkh);
  
  not rkduoajguu(qb, oitb);
  
  or azju(nfxlbumnpw, yjzbzu, eovcuyo);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint eovcuyo -> logic eovcuyo
  
  
  // Single-driven assigns
  assign mrcyxwzl = '{'{'{'b00111}},'{'{'b01001}},'{'{'b10000}},'{'{'b1100}}};
  assign lns = lns;
  
  // Multi-driven assigns
  assign yjzbzu = eovcuyo;
  assign oitb = oitb;
  assign syferkh = 'b1;
  assign hbfehdouq = eovcuyo;
endmodule: wvmtb

module bvwsab
  (output longint eqoh);
  
  
  not ayaf(wji, nekhxtuox);
  
  xor wrx(ni, o, eqoh);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint eqoh -> logic eqoh
  
  not lfezlr(o, ni);
  
  xor gvrsvpa(nekhxtuox, ni, nekhxtuox);
  
  
  // Single-driven assigns
  assign eqoh = nekhxtuox;
  
  // Multi-driven assigns
  assign o = 'b1;
  assign ni = nekhxtuox;
  assign wji = eqoh;
endmodule: bvwsab



// Seed after: 12658144569597683733,3128299129089410139
