// Seed: 9931058363952773939,3128299129089410139

module w
  (output reg biryrjfbif [1:1], output logic [1:4] skmdql [3:2][0:2][2:2], output wand logic [1:0][2:1][2:3][1:3] g [0:1][3:3][2:4]);
  
  
  not nzxt(rt, r);
  
  or xlqx(vdawvpw, r, opxaf);
  
  xor furqxtq(dwhgohg, kypkpr, dwhgohg);
  
  xor koghkulf(r, r, ifqjhz);
  
  
  // Single-driven assigns
  assign skmdql = '{'{'{'{'b11zzx,'bx10z,'b101x,'bxxzx0}},'{'{'b1011,'bx,'b0z100,'bzz0}},'{'{'b111,'b1z0z,'bx0x,'b1}}},'{'{'{'b01xz1,'b1x00,'b1x,'bx1}},'{'{'bx00x,'bxz0z,'bxzx,'b10x}},'{'{'b0,'bxxxx,'b1x1xz,'b01z1z}}}};
  assign biryrjfbif = biryrjfbif;
  
  // Multi-driven assigns
  assign g = g;
  assign opxaf = 'b0;
  assign r = 'b0;
  assign vdawvpw = 'bxz0x;
  assign ifqjhz = rt;
endmodule: w

module vqhoakr
  (output reg [3:0] a [0:1], output logic [4:0][0:1][2:1][3:0]  uht, output time ytniovkvde [0:0], output time n);
  
  
  not mo(uht, wfe);
  // warning: implicit conversion of port connection expands from 1 to 80 bits
  //   logic uht -> logic [4:0][0:1][2:1][3:0]  uht
  
  not mnmfuo(mtycpdq, ctusm);
  
  or aqcml(n, jlzvfbfb, tiynzcbvvm);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  //   logic n -> time n
  
  
  // Single-driven assigns
  assign a = a;
  assign ytniovkvde = '{'b1x0z};
  
  // Multi-driven assigns
  assign wfe = 'bx100;
  assign tiynzcbvvm = 'bx;
  assign ctusm = 'b0;
endmodule: vqhoakr

module vbfuvlwh
  ( output tri logic [3:0][4:4][2:4] dstlzlj [4:4][2:2][4:4]
  , input wire logic [3:4][1:1] en [0:4][0:4][2:1][3:3]
  , input bit [2:3][2:3][3:1]  qicozo
  , input logic [0:2][2:1] zbgcveaku [3:3][0:0]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign en = en;
  assign dstlzlj = dstlzlj;
endmodule: vbfuvlwh



// Seed after: 4773139017576541913,3128299129089410139
