// Seed: 2775971243336691657,3128299129089410139

module ty
  ( output logic olplrepxh [1:1]
  , output trior logic [2:0][4:3][0:3][1:0] vdd [2:4][4:3][2:0][2:4]
  , input wire logic yimanrlpqz
  , input logic [0:1][4:2][0:2]  skhkqzigv
  , input bit qweuypel [2:2]
  , input reg [0:4][0:1]  xb
  );
  
  
  or sjt(gc, yimanrlpqz, yimanrlpqz);
  
  not jzyncfbwm(yimanrlpqz, skhkqzigv);
  // warning: implicit conversion of port connection truncates from 18 to 1 bits
  //   logic [0:1][4:2][0:2]  skhkqzigv -> logic skhkqzigv
  
  xor bmqhclkti(yimanrlpqz, yimanrlpqz, yimanrlpqz);
  
  or efsm(gxmzank, xb, gc);
  // warning: implicit conversion of port connection truncates from 10 to 1 bits
  //   reg [0:4][0:1]  xb -> logic xb
  
  
  // Single-driven assigns
  assign olplrepxh = '{'bzz0};
  
  // Multi-driven assigns
  assign vdd = vdd;
  assign gc = 'bx;
  assign yimanrlpqz = 'bz;
  assign gxmzank = xb;
endmodule: ty

module lrjsagnzj
  ( output uwire logic [4:1][1:1][1:0] aophfxii [0:0][1:4][1:2][0:3]
  , output bit enfi
  , input tri1 logic [3:3][2:3][0:3] ihh [1:3][0:1][1:0]
  , input supply1 logic q [0:3]
  );
  
  
  not hpsiip(kr, vorflsd);
  
  nand h(enfi, enfi, enfi);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic enfi -> bit enfi
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit enfi -> logic enfi
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit enfi -> logic enfi
  
  nand ewmhx(vorflsd, vorflsd, enfi);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit enfi -> logic enfi
  
  
  // Single-driven assigns
  assign aophfxii = aophfxii;
  
  // Multi-driven assigns
endmodule: lrjsagnzj

module glnxp
  (output tri0 logic [3:2] ervhu [2:3][4:2], input reg [3:3][2:3] fnr [4:3][4:0], input wire logic [0:1]  en, input logic [1:0]  y);
  
  
  or jea(debwxgxugl, debwxgxugl, debwxgxugl);
  
  not obvvkzvp(rdnrjyd, debwxgxugl);
  
  and nuqz(debwxgxugl, vbgnryz, oymxownm);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ervhu = ervhu;
  assign vbgnryz = en;
endmodule: glnxp

module wubhfsqb
  (output tri1 logic [0:3][1:2] ge [0:4][2:3][0:0], input logic nweae [2:2]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ge = ge;
endmodule: wubhfsqb



// Seed after: 1772075317299193651,3128299129089410139
