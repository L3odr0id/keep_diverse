// Seed: 13160880725827085634,3128299129089410139

module vxhilwa
  ( output wire logic [4:3][4:4][1:2] uagcy [3:2][3:4][3:3]
  , output reg [3:3] kbzgyzrrti [0:0]
  , output reg [1:4][1:3][4:3][3:2]  ix
  , output logic [3:2][3:3][2:0][0:3]  axkgemuj
  , input tri0 logic [0:2][4:0][0:1][1:1] olmboy [3:4][4:1][4:4]
  , input logic mnm
  );
  
  
  
  // Single-driven assigns
  assign kbzgyzrrti = '{'{'bx1z}};
  assign ix = '{'{'{'{'b0,'b1},'{'bx0x1,'bxz1}},'{'{'bx1,'bx},'{'b1z0,'b0zz}},'{'{'b0,'b11xx},'{'bxxxz,'bxxxx}}},'{'{'{'b0,'bxz10},'{'bz01z0,'bzz0}},'{'{'bx1zz1,'b1xx10},'{'bz1zx,'bx0xx}},'{'{'b0zzz,'b1},'{'b01x,'b0xzz}}},'{'{'{'b100xx,'b0},'{'bx,'bx11x0}},'{'{'b11,'bx01},'{'bz,'bz0zx}},'{'{'b101,'b0},'{'b1z011,'bxz1}}},'{'{'{'bz0zz0,'bz},'{'bzx,'b0x1x1}},'{'{'bz11xz,'b11},'{'b00z1,'bx0010}},'{'{'b00x1x,'b0xz0z},'{'bzx,'b0x0x1}}}};
  assign axkgemuj = '{'{'{'{'b1,'bx0zxx,'b0z,'b1},'{'bz,'b1xx1x,'bx1z,'bx1xx},'{'b00zzx,'b0xz1,'b00z1,'bz}}},'{'{'{'b01,'bz11z1,'bz,'b111xz},'{'b1x10x,'bzx010,'b1x,'bx},'{'bx1,'b0,'b100xx,'b0z}}}};
  
  // Multi-driven assigns
endmodule: vxhilwa

module hnzkccny
  (output tri logic [0:1][0:1]  rdxvxksh, output reg [0:1][1:4][3:2]  aqwu);
  
  
  not pu(rdxvxksh, aqwu);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic rdxvxksh -> tri logic [0:1][0:1]  rdxvxksh
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   reg [0:1][1:4][3:2]  aqwu -> logic aqwu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rdxvxksh = rdxvxksh;
endmodule: hnzkccny



// Seed after: 8128931952326600637,3128299129089410139
