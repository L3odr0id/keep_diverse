// Seed: 4919911431090630944,3128299129089410139

module y
  ( output uwire logic [1:2][0:1][0:0][1:0] okgqrdn [0:1][4:3][2:1]
  , output reg iwvnjkmjx
  , output tri0 logic [0:3][3:0][4:1]  rtoher
  , input bit [4:1][4:2][2:2]  skcmhwk
  , input uwire logic [0:1]  savw
  , input logic [3:1]  yjzn
  );
  
  
  and smjyv(izgexfhs, savw, iwvnjkmjx);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   uwire logic [0:1]  savw -> logic savw
  
  
  // Single-driven assigns
  assign okgqrdn = okgqrdn;
  assign iwvnjkmjx = iwvnjkmjx;
  
  // Multi-driven assigns
  assign izgexfhs = 'b0x000;
  assign rtoher = iwvnjkmjx;
endmodule: y

module gvpkmfe
  ( output byte cgdkcqogd [4:2]
  , output wor logic [1:3][4:1] kjgmmxavd [3:4][1:4][1:4]
  , output trireg logic [4:1][3:2][3:0][0:1] jzohsgncvh [3:4][2:1][4:0]
  , input logic [0:4] fqsvezuk [0:4]
  , input triand logic [3:4][1:1][3:0][0:0]  jjaybu
  , input tri0 logic [0:0][3:3][3:3] srdset [4:2]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jzohsgncvh = jzohsgncvh;
  assign jjaybu = '{'{'{'{'b0z},'{'bzz1},'{'b00z0},'{'b01}}},'{'{'{'b1xz0},'{'bx00x},'{'b11},'{'b0}}}};
  assign kjgmmxavd = kjgmmxavd;
  assign srdset = srdset;
endmodule: gvpkmfe



// Seed after: 7084504391126471160,3128299129089410139
