// Seed: 2769780858164702270,3128299129089410139

module df
  (output triand logic [3:3] doasrorij [4:0][1:1], input reg [0:2][2:1]  zfhourck, input wand logic [4:0]  dr);
  
  
  not npriepkaa(payw, dr);
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   wand logic [4:0]  dr -> logic dr
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign doasrorij = '{'{'{'b0}},'{'{'bxzxz}},'{'{'b1x0}},'{'{'b1xx}},'{'{'b1x}}};
  assign dr = dr;
endmodule: df

module mehhebl
  (output trior logic [0:4][2:3] ghsv [4:1][1:3]);
  
  triand logic [3:3] bdljzxyyhu [4:0][1:1];
  
  or rpscmct(igv, wwop, wwop);
  
  not bm(ttmxlxaaui, r);
  
  not u(igv, r);
  
  df uvafsa(.doasrorij(bdljzxyyhu), .zfhourck(xuczggn), .dr(wwop));
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   wire logic xuczggn -> reg [0:2][2:1]  zfhourck
  //
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   wire logic wwop -> wand logic [4:0]  dr
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ghsv = '{'{'{'{'bxz100,'bxx},'{'b0zxx,'bxxz00},'{'bz1001,'b1x01},'{'bxx1x,'bx},'{'b0,'b00}},'{'{'b10x,'bz01},'{'bx101x,'bz},'{'b1,'bzzx},'{'b0z1z,'bx},'{'bz1,'b0}},'{'{'bx1zz0,'b00},'{'b11zx,'b1zz10},'{'b0,'bz},'{'bz,'b1},'{'b1,'b00}}},'{'{'{'bz10,'bxz1xx},'{'bx01x,'b01110},'{'bzx,'bzz1xx},'{'b01x0,'bzx},'{'b10z1,'b1z00}},'{'{'b0zxxz,'bxz0z0},'{'b0z,'bz1111},'{'b0zx,'b0100},'{'b1x,'b1zx1},'{'bzz,'b0zx}},'{'{'b1010,'bz0},'{'bxx,'b011x},'{'bx,'b10x},'{'b10z,'bzzx0},'{'b1z,'bxz010}}},'{'{'{'bx11,'b0z0},'{'bxzx01,'bx0xx},'{'bz11z,'b01},'{'b110x,'bx},'{'b1,'bzx0}},'{'{'bz1x,'bz1},'{'b0z1z,'bz},'{'b100xx,'b0xx},'{'b0z1,'bxxx},'{'b00,'bz}},'{'{'b1xxz1,'bzxxxz},'{'b0x00,'bxz},'{'b1,'bx0xz},'{'bzx11,'bxz11},'{'b01zz,'bzzzx0}}},'{'{'{'b0,'b1},'{'bzx0,'b0x},'{'b0xx1z,'bz},'{'b00,'b1xzz},'{'bx,'bz}},'{'{'b1zx1,'bx100},'{'b0x0z,'bz1z0},'{'bxz11,'bz0xx},'{'b0,'b1x},'{'b01z1z,'b1x}},'{'{'bx01z1,'bx},'{'b1x00z,'b1z},'{'b1zzxx,'b1z},'{'bz,'b0},'{'bz010,'bz110}}}};
  assign xuczggn = 'bx0z;
  assign r = wwop;
  assign wwop = xuczggn;
endmodule: mehhebl

module czwp
  (input triand logic [0:3][2:0][1:2][1:2]  wh);
  
  triand logic [3:3] og [4:0][1:1];
  triand logic [3:3] zonq [4:0][1:1];
  
  df ntydsrfjxp(.doasrorij(zonq), .zfhourck(wh), .dr(orwqo));
  // warning: implicit conversion of port connection truncates from 48 to 6 bits
  //   triand logic [0:3][2:0][1:2][1:2]  wh -> reg [0:2][2:1]  zfhourck
  //
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   wire logic orwqo -> wand logic [4:0]  dr
  
  and dvne(wh, wh, wh);
  // warning: implicit conversion of port connection expands from 1 to 48 bits
  //   logic wh -> triand logic [0:3][2:0][1:2][1:2]  wh
  //
  // warning: implicit conversion of port connection truncates from 48 to 1 bits
  //   triand logic [0:3][2:0][1:2][1:2]  wh -> logic wh
  //
  // warning: implicit conversion of port connection truncates from 48 to 1 bits
  //   triand logic [0:3][2:0][1:2][1:2]  wh -> logic wh
  
  df cuy(.doasrorij(og), .zfhourck(zzq), .dr(kirgoye));
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   wire logic zzq -> reg [0:2][2:1]  zfhourck
  //
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   wire logic kirgoye -> wand logic [4:0]  dr
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign orwqo = 'b000;
endmodule: czwp

module ahoyjk
  ( output supply0 logic [3:2][4:2][1:0] dwj [0:4]
  , output wire logic [1:0][2:4] thrkcwpqo [0:2][2:4][3:0][0:3]
  , input wor logic [0:2] lmx [4:3][3:0][3:4][2:4]
  );
  
  
  not ieq(lvjdi, lvjdi);
  
  not fwtjch(lvjdi, lvjdi);
  
  not mnbz(lvjdi, jxtasmng);
  
  and pjr(lvjdi, lvjdi, lvjdi);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dwj = dwj;
endmodule: ahoyjk



// Seed after: 11800529220501756588,3128299129089410139
