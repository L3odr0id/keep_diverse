// Seed: 8699459758548135104,3128299129089410139

module ewfhqxg
  ( output time vbpt
  , output reg [0:0][2:4][0:1][3:4]  ebvsol
  , output tri0 logic dligbsq [3:4][3:2][2:4]
  , input tri1 logic dawpxivzdi [1:0][3:1][1:2]
  , input uwire logic [1:4] vqtgqlcm [0:1][4:0]
  , input trireg logic [2:0][3:4][4:1] tkfnakrg [0:4]
  );
  
  
  or wm(tlwpbkvvsv, tlwpbkvvsv, ebvsol);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [0:0][2:4][0:1][3:4]  ebvsol -> logic ebvsol
  
  or biwb(ezax, vbpt, sqjhkem);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time vbpt -> logic vbpt
  
  nand fabmcmez(kuejxglrra, w, qplp);
  
  or ebcoealak(v, vterjlia, v);
  
  
  // Single-driven assigns
  assign vbpt = vbpt;
  assign ebvsol = qplp;
  
  // Multi-driven assigns
endmodule: ewfhqxg



// Seed after: 15337481340297115087,3128299129089410139
