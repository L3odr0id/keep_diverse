// Seed: 3035589897675090996,3128299129089410139

module tcnwioc
  ( output triand logic [3:4][2:4] hgyenq [1:3][1:2]
  , input time loddtn [0:2][0:4]
  , input reg [2:3][0:2][2:4][2:0]  uzneel
  , input reg [1:1][2:2]  gvgsqe
  , input triand logic [1:0] eiolcbjq [2:3][2:4][3:2][2:0]
  );
  
  
  or ntpnkhtnc(gyzcfxxik, uzneel, gvgsqe);
  // warning: implicit conversion of port connection truncates from 54 to 1 bits
  //   reg [2:3][0:2][2:4][2:0]  uzneel -> logic uzneel
  
  not sdqjzqbvwg(inifolp, gyzcfxxik);
  
  nand dn(hmdcsrizh, hq, uzneel);
  // warning: implicit conversion of port connection truncates from 54 to 1 bits
  //   reg [2:3][0:2][2:4][2:0]  uzneel -> logic uzneel
  
  not mtni(lux, hmdcsrizh);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hgyenq = hgyenq;
  assign eiolcbjq = eiolcbjq;
  assign hq = 'b1z01;
  assign hmdcsrizh = gvgsqe;
  assign gyzcfxxik = uzneel;
endmodule: tcnwioc



// Seed after: 14973839198957523227,3128299129089410139
