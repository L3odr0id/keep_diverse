// Seed: 16560062601981626402,3128299129089410139

module uyb
  (input reg [4:4][0:2]  nptxaarju, input supply0 logic [2:0][0:0][3:1][1:4] fm [2:4], input logic [4:0][2:1] dxqfe [0:3]);
  
  
  not tvw(jershq, q);
  
  or hsqyvv(ccfrf, ccfrf, q);
  
  xor sapud(q, ccfrf, nptxaarju);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [4:4][0:2]  nptxaarju -> logic nptxaarju
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign q = 'bz1;
  assign jershq = ccfrf;
  assign fm = fm;
  assign ccfrf = q;
endmodule: uyb

module zunqizydu
  ( output shortint dtfjyjfo [1:2][3:4]
  , output wor logic [1:2]  uxhhv
  , output longint u
  , input triand logic [3:2] nbxowrj [4:4][4:1]
  , input tri logic yc [3:1][0:4][2:3]
  , input trior logic [0:3][0:2][4:0][0:0] i [3:4][4:0]
  );
  
  
  and qqyl(uxhhv, uxhhv, uxhhv);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic uxhhv -> wor logic [1:2]  uxhhv
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   wor logic [1:2]  uxhhv -> logic uxhhv
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   wor logic [1:2]  uxhhv -> logic uxhhv
  
  
  // Single-driven assigns
  assign dtfjyjfo = '{'{'b01,'b011},'{'b0111,'b1}};
  assign u = uxhhv;
  
  // Multi-driven assigns
  assign uxhhv = '{'b0,'bxx};
endmodule: zunqizydu



// Seed after: 10701314730660828924,3128299129089410139
