// Seed: 11378901856138186289,3128299129089410139

module b
  ( output reg [4:3]  bhi
  , output byte hfxcn
  , input logic [0:3]  tspathqrnb
  , input tri0 logic [4:1][4:3][1:2]  hnzhkipil
  , input logic [1:4][4:0][3:0][3:1]  txood
  , input wand logic [1:1][4:3] zfzhfayppj [2:1]
  );
  
  
  and mddw(ibpz, hnzhkipil, txood);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   tri0 logic [4:1][4:3][1:2]  hnzhkipil -> logic hnzhkipil
  //
  // warning: implicit conversion of port connection truncates from 240 to 1 bits
  //   logic [1:4][4:0][3:0][3:1]  txood -> logic txood
  
  not n(yxvizxmdy, bhi);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   reg [4:3]  bhi -> logic bhi
  
  or vstass(utirkxqb, hpjxqyce, iu);
  
  and tacnrnyck(cykrzaowvt, ypssool, biiy);
  
  
  // Single-driven assigns
  assign bhi = bhi;
  assign hfxcn = 'b0110;
  
  // Multi-driven assigns
  assign utirkxqb = utirkxqb;
  assign ibpz = hnzhkipil;
  assign yxvizxmdy = 'bzzxz1;
  assign hnzhkipil = hnzhkipil;
  assign zfzhfayppj = '{'{'{'b01z,'b1zx}},'{'{'b0,'b00xx}}};
endmodule: b

module m
  ( output tri logic [0:0][3:4] hcmsfue [3:1][1:1][2:3]
  , output trior logic [3:2][2:3] oea [0:0][2:4]
  , output logic [4:3][4:0]  hbmuyo
  , output reg [0:1][0:1][4:0] gimodgc [4:4]
  , input tri1 logic [3:3] mxrlgtqvd [4:1][4:1][4:0][0:1]
  , input tri logic [0:3][1:0] hcepwddzmp [0:4][4:2]
  );
  
  
  
  // Single-driven assigns
  assign hbmuyo = hbmuyo;
  assign gimodgc = '{'{'{'{'b11,'b01x,'b11,'b1,'bz1x},'{'bxz00x,'bx1z0,'bzxzz1,'bx01x,'b0}},'{'{'bx00z,'bx0zxz,'bxx10z,'b00,'bx},'{'bzzxx,'bz00,'b1x10,'b1zxz,'b11100}}}};
  
  // Multi-driven assigns
  assign hcepwddzmp = hcepwddzmp;
endmodule: m



// Seed after: 4868562018233217693,3128299129089410139
