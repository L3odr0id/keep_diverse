// Seed: 5245149075574092761,3128299129089410139

module ihhh
  (output tri logic [4:2][2:2][3:2][2:0] kvd [2:4]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kvd = kvd;
endmodule: ihhh

module kgxhpjb
  ();
  
  
  xor lpvxqkatd(mzgshbhu, eu, eu);
  
  not mvqlumhcy(eu, eu);
  
  not dway(xqt, zg);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign eu = zg;
  assign zg = mzgshbhu;
  assign mzgshbhu = zg;
endmodule: kgxhpjb

module wfomqgdtx
  ( output wire logic [1:3] uikn [3:2][0:1][4:3][4:0]
  , output logic [0:1][4:4][3:4]  febhrckma
  , output bit ojj
  , input triand logic l [0:1][0:1]
  , input integer dwxulilk [2:2]
  );
  
  
  nand a(no, febhrckma, on);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   logic [0:1][4:4][3:4]  febhrckma -> logic febhrckma
  
  
  // Single-driven assigns
  assign ojj = 'b1110;
  assign febhrckma = '{'{'{'b01x0z,'b011}},'{'{'bx,'b1xxx0}}};
  
  // Multi-driven assigns
endmodule: wfomqgdtx



// Seed after: 16610296227259165878,3128299129089410139
