// Seed: 1772075317299193651,3128299129089410139

module tqz
  ( output uwire logic [2:2][2:3][4:3] faulofgbok [4:0][1:1][4:4][3:1]
  , input trireg logic [1:2][1:2][3:0][1:0] shvugfvt [4:0][1:1][0:3][4:1]
  , input reg [1:1][3:0][3:3][3:0]  bo
  );
  
  
  nand brxuze(ejwnnvenu, ejwnnvenu, usnztvbah);
  
  not ethzf(usnztvbah, usnztvbah);
  
  and qmltcwzmv(kjf, txmxb, dwrglchkug);
  
  
  // Single-driven assigns
  assign faulofgbok = faulofgbok;
  
  // Multi-driven assigns
  assign ejwnnvenu = 'bz0;
endmodule: tqz

module daccsinzk
  (output trior logic [4:2]  sma, output logic [0:2][2:0][4:0][2:2]  u, output tri1 logic ziqo [4:4][4:0][3:4]);
  
  
  not sue(mzha, blqgaftn);
  
  
  // Single-driven assigns
  assign u = u;
  
  // Multi-driven assigns
  assign sma = u;
  assign mzha = sma;
  assign blqgaftn = sma;
  assign ziqo = ziqo;
endmodule: daccsinzk

module oxo
  ( output shortint tnlwybac [1:0]
  , output bit [0:4] qg [0:0][4:0][2:1]
  , input uwire logic [0:2][1:1][4:0] ai [3:2]
  , input logic [1:4][3:2][3:1]  rhd
  );
  
  
  not fnbzaktwm(lo, rhd);
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   logic [1:4][3:2][3:1]  rhd -> logic rhd
  
  
  // Single-driven assigns
  assign qg = qg;
  assign tnlwybac = tnlwybac;
  
  // Multi-driven assigns
  assign lo = 'bxx;
endmodule: oxo



// Seed after: 9099988925635228673,3128299129089410139
