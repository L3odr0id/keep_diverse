// Seed: 15923648016595859751,3128299129089410139

module oi
  ( output uwire logic iilbvakv [4:2]
  , output bit [3:3][1:1]  lw
  , output uwire logic [3:2] cd [4:2][0:3][1:0]
  , input wor logic [2:0][2:0][3:2] kpjijejdr [0:2]
  , input trior logic [0:1][2:2] rlgx [0:0][4:3][3:3][3:2]
  , input realtime vlkzlivo [3:1][1:1]
  );
  
  
  not cixjvmoctm(lw, lw);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic lw -> bit [3:3][1:1]  lw
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:3][1:1]  lw -> logic lw
  
  and xp(syi, lw, zjmw);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:3][1:1]  lw -> logic lw
  
  
  // Single-driven assigns
  assign cd = cd;
  assign iilbvakv = '{'bx0z10,'bzxz00,'bx0z};
  
  // Multi-driven assigns
  assign zjmw = 'bz001z;
  assign syi = lw;
  assign rlgx = rlgx;
  assign kpjijejdr = kpjijejdr;
endmodule: oi

module npchnew
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: npchnew

module pweaqa
  ( output tri logic [0:0][2:1] uq [3:3][0:2]
  , input tri logic ji [2:4][2:0][1:3][1:1]
  , input tri logic [0:4][3:1][0:1][0:0] nmvseoe [1:2][2:1][1:2][2:4]
  , input bit [2:2] a [2:1][0:2]
  , input logic hroizuxt [4:4][4:3][2:1]
  );
  
  
  and lc(prraxaivbb, casysgglob, qvpmorlbly);
  
  or nwgc(kqkidrta, hkekmh, ailaf);
  
  xor rc(prraxaivbb, wv, ufcfnvyf);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: pweaqa



// Seed after: 16013029700436987217,3128299129089410139
