// Seed: 12822400028629458463,3128299129089410139

module w
  ( output wor logic [0:2]  hhgljaumo
  , input bit [3:0][1:1][0:0]  hnxlb
  , input triand logic [1:3][1:0][1:1] svzqqr [4:3][2:4][1:1][0:4]
  , input reg [1:0]  lgaplwcqvh
  , input triand logic [0:0][2:2][0:4] rbvhjkwt [2:3][3:0][1:3][3:2]
  );
  
  
  and dkaemsber(hhgljaumo, hhgljaumo, hhgljaumo);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic hhgljaumo -> wor logic [0:2]  hhgljaumo
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wor logic [0:2]  hhgljaumo -> logic hhgljaumo
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wor logic [0:2]  hhgljaumo -> logic hhgljaumo
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hhgljaumo = '{'b1xz1,'bx,'bzzxz};
endmodule: w

module kydjqm
  (output shortint wjpjug, output logic wwgye, input logic [2:0][2:1][2:4][0:1]  l);
  
  
  and kj(wwgye, wjpjug, l);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint wjpjug -> logic wjpjug
  //
  // warning: implicit conversion of port connection truncates from 36 to 1 bits
  //   logic [2:0][2:1][2:4][0:1]  l -> logic l
  
  not hgd(wjpjug, nr);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic wjpjug -> shortint wjpjug
  
  and tg(annrtuffk, sbzslse, wwgye);
  
  not aa(khou, l);
  // warning: implicit conversion of port connection truncates from 36 to 1 bits
  //   logic [2:0][2:1][2:4][0:1]  l -> logic l
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nr = 'b0;
  assign annrtuffk = 'bzxx;
  assign khou = wjpjug;
  assign sbzslse = wjpjug;
endmodule: kydjqm



// Seed after: 16536538239648392389,3128299129089410139
