// Seed: 7075531678909538591,3128299129089410139

module bulos
  ( output wand logic znwdyroq
  , output tri1 logic dspkb [2:4][2:4][3:1]
  , output trireg logic [0:1][0:4] wrqyydhc [4:1][2:3][3:1]
  , output bit [3:2][1:2]  kfmtafnek
  , input realtime nrtvod
  , input tri logic [1:4][2:3] tbpljjuybe [0:0]
  , input uwire logic [2:3][3:3][0:1] hyvobzjirw [2:0][0:2]
  , input tri0 logic [2:2] gs [2:0][1:0][1:2]
  );
  
  
  xor acadh(epqscfp, ickfpiuu, znwdyroq);
  
  
  // Single-driven assigns
  assign kfmtafnek = epqscfp;
  
  // Multi-driven assigns
endmodule: bulos



// Seed after: 574283273884231197,3128299129089410139
