// Seed: 5555284318056057502,3128299129089410139

module ak
  (output real vfcbx [4:2][1:4][2:3], output bit veh [2:3][2:2], output bit [3:4][4:1] xnpvgjgwm [4:3]);
  
  
  and alljf(bioza, bioza, aghjfwnyf);
  
  
  // Single-driven assigns
  assign vfcbx = '{'{'{'b1,'bz},'{'bxxxz0,'b1},'{'b011z,'bx111},'{'bxzz0,'bzz1x}},'{'{'b1010z,'b0z},'{'bx11z,'b00z},'{'b1xzxz,'b0101},'{'bz1z0,'b1xx}},'{'{'b1z,'bxzz},'{'b1,'bxz00},'{'bzzzz,'bxz1z0},'{'bxz0,'bzz1}}};
  assign veh = '{'{'b0101},'{'b10111}};
  
  // Multi-driven assigns
  assign aghjfwnyf = 'b000;
  assign bioza = 'b01x1;
endmodule: ak

module bkf
  ( input wire logic [4:1][4:0][4:1] zhn [0:0][1:0][2:1][0:1]
  , input shortreal jreqjj
  , input bit [3:4] hddils [1:2]
  , input bit [0:2][1:0][1:1][0:0]  rdjsjhqatr
  );
  
  
  not ijvq(lo, cuc);
  
  or ixdaytgk(zuxqoj, cuc, xvmrzbad);
  
  nand u(cuc, sew, sew);
  
  not bbenjc(cuc, cuc);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zhn = zhn;
  assign sew = cuc;
  assign xvmrzbad = 'bz;
  assign cuc = 'b0x000;
endmodule: bkf

module qadyerc
  (output bit [3:0][3:3]  h, input tri logic [0:4][0:1]  tga, input bit [1:2][1:3][0:0]  ztvmhdj, input real node);
  
  bit [3:4] wohlwfg [1:2];
  wire logic [4:1][4:0][4:1] oikfhifxu [0:0][1:0][2:1][0:1];
  
  not mdgml(tga, h);
  // warning: implicit conversion of port connection expands from 1 to 10 bits
  //   logic tga -> tri logic [0:4][0:1]  tga
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:0][3:3]  h -> logic h
  
  bkf saknvqex(.zhn(oikfhifxu), .jreqjj(h), .hddils(wohlwfg), .rdjsjhqatr(h));
  // warning: implicit conversion of port connection expands from 4 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:0][3:3]  h -> shortreal jreqjj
  //
  // warning: implicit conversion of port connection expands from 4 to 6 bits
  //   bit [3:0][3:3]  h -> bit [0:2][1:0][1:1][0:0]  rdjsjhqatr
  
  
  // Single-driven assigns
  assign wohlwfg = '{'{'b010,'b110},'{'b0,'b00}};
  
  // Multi-driven assigns
  assign oikfhifxu = oikfhifxu;
endmodule: qadyerc

module ha
  (input bit [4:1][1:0] qqajakupjd [0:4][2:0], input logic [1:1][2:1] geygj [1:2][1:3]);
  
  bit [3:4][4:1] ww [4:3];
  bit u [2:3][2:2];
  real cqur [4:2][1:4][2:3];
  
  ak dquaifizy(.vfcbx(cqur), .veh(u), .xnpvgjgwm(ww));
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ha



// Seed after: 4261191817767376468,3128299129089410139
