// Seed: 11691253499933042360,3128299129089410139

module rggtow
  ( output logic [4:1][1:1][4:1][4:0]  uyxmdp
  , input bit [4:4] kpp [4:0]
  , input supply0 logic [2:2][0:3][2:3] rqtyhdu [4:2][1:1][4:3][1:2]
  );
  
  
  nand jqtxgts(ijzegsab, ijzegsab, khthwpyg);
  
  not rqtebdt(ijzegsab, oswdp);
  
  not ashz(ijzegsab, uyxmdp);
  // warning: implicit conversion of port connection truncates from 80 to 1 bits
  //   logic [4:1][1:1][4:1][4:0]  uyxmdp -> logic uyxmdp
  
  not c(fmqlfcatrl, kyilybcwu);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: rggtow

module gpr
  (output shortint j [1:4]);
  
  
  not avd(gmd, muxfijc);
  
  not ityjj(gmd, muxfijc);
  
  nand jxes(gmd, muxfijc, muxfijc);
  
  
  // Single-driven assigns
  assign j = '{'b0001,'b10100,'b010,'b00000};
  
  // Multi-driven assigns
  assign gmd = 'b0x;
  assign muxfijc = 'b1zz1x;
endmodule: gpr

module nayunfph
  (output logic [1:3][4:2] zwaptqlzw [2:4], output shortreal iwh, output triand logic clrrm [1:3][0:0], input bit jvblg);
  
  
  not uty(iwh, r);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic iwh -> shortreal iwh
  
  
  // Single-driven assigns
  assign zwaptqlzw = zwaptqlzw;
  
  // Multi-driven assigns
  assign clrrm = clrrm;
endmodule: nayunfph



// Seed after: 13510878130923757581,3128299129089410139
