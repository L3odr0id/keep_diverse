// Seed: 2189224357496412630,3128299129089410139

module zswzjadvn
  (output tri logic [0:4][2:3][3:0] h [0:1][0:1][4:1], output supply0 logic [1:1][4:0][4:1][1:0]  qygsew);
  
  
  not sio(qygsew, qygsew);
  // warning: implicit conversion of port connection expands from 1 to 40 bits
  //   logic qygsew -> supply0 logic [1:1][4:0][4:1][1:0]  qygsew
  //
  // warning: implicit conversion of port connection truncates from 40 to 1 bits
  //   supply0 logic [1:1][4:0][4:1][1:0]  qygsew -> logic qygsew
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign h = h;
  assign qygsew = '{'{'{'{'bz0x1,'bx1000},'{'bxx011,'b111xx},'{'bz0x,'bz10},'{'bz0z0,'bzz0z}},'{'{'bzzz,'b1},'{'b1xzzx,'bx10xx},'{'bzx,'bx},'{'bxx,'b0x0z}},'{'{'b0,'b0xx1z},'{'bxz,'bx10},'{'bz0xz,'b10},'{'b11z,'b00xx}},'{'{'b0,'b1zzxz},'{'bx1z,'b11},'{'b1,'bz},'{'bzx10,'b0}},'{'{'b0x,'b1zz0},'{'b00,'b00xx},'{'b0z1,'bzz0x1},'{'bzz,'bz}}}};
endmodule: zswzjadvn

module w
  ( output wor logic [4:1][0:2][4:0]  e
  , output bit [4:0]  jsot
  , output trior logic [3:2][3:4][1:4]  dkcfaui
  , input byte sxwo
  , input wire logic [3:1] vura [0:2][2:1][3:0][3:1]
  , input supply1 logic [3:2] rhcowfqs [0:1][3:4][0:0]
  );
  
  tri logic [0:4][2:3][3:0] zgtvgs [0:1][0:1][4:1];
  
  zswzjadvn rhm(.h(zgtvgs), .qygsew(renr));
  // warning: implicit conversion of port connection truncates from 40 to 1 bits
  //   supply0 logic [1:1][4:0][4:1][1:0]  qygsew -> wire logic renr
  
  not rb(svagpu, dh);
  
  or bsav(e, e, fg);
  // warning: implicit conversion of port connection expands from 1 to 60 bits
  //   logic e -> wor logic [4:1][0:2][4:0]  e
  //
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   wor logic [4:1][0:2][4:0]  e -> logic e
  
  nand gyit(wajkohz, dj, imlsbb);
  
  
  // Single-driven assigns
  assign jsot = e;
  
  // Multi-driven assigns
  assign zgtvgs = zgtvgs;
  assign dj = 'b00z;
endmodule: w

module ixi
  ( output logic [3:0][3:4][1:1]  lt
  , output tri logic [4:0][4:3][3:0][3:1] qbu [2:4]
  , input time vclllhbuuh
  , input logic [1:3][2:4][1:3][2:4]  pgzvid
  , input supply0 logic [1:1][2:0][3:4][3:1] ataym [1:4][4:4][4:4]
  , input reg [2:2][1:3][2:3]  kdyziobqu
  );
  
  supply1 logic [3:2] ce [0:1][3:4][0:0];
  wire logic [3:1] onzbkikzle [0:2][2:1][3:0][3:1];
  
  not mylggpkwhe(lt, lt);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   logic lt -> logic [3:0][3:4][1:1]  lt
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   logic [3:0][3:4][1:1]  lt -> logic lt
  
  nand uxxqvtrt(poqmmzy, lt, pgzvid);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   logic [3:0][3:4][1:1]  lt -> logic lt
  //
  // warning: implicit conversion of port connection truncates from 81 to 1 bits
  //   logic [1:3][2:4][1:3][2:4]  pgzvid -> logic pgzvid
  
  w uwjom(.e(wqqdkf), .jsot(dcrskeiixy), .dkcfaui(sgjbntxzch), .sxwo(pgzvid), .vura(onzbkikzle), .rhcowfqs(ce));
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   wor logic [4:1][0:2][4:0]  e -> wire logic wqqdkf
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:0]  jsot -> wire logic dcrskeiixy
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   trior logic [3:2][3:4][1:4]  dkcfaui -> wire logic sgjbntxzch
  //
  // warning: implicit conversion of port connection truncates from 81 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic [1:3][2:4][1:3][2:4]  pgzvid -> byte sxwo
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign sgjbntxzch = lt;
  assign qbu = qbu;
  assign dcrskeiixy = lt;
endmodule: ixi



// Seed after: 12822400028629458463,3128299129089410139
