// Seed: 16755045049282625894,3128299129089410139

module mf
  ( input logic [1:4] t [0:2][3:0][1:2]
  , input realtime qthncx
  , input triand logic [4:3][4:2][1:0][0:4]  xxptc
  , input wire logic vwsbam [1:4][4:0][1:0][3:2]
  );
  
  
  not lc(wz, qthncx);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime qthncx -> logic qthncx
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign wz = 'bz0;
  assign xxptc = '{'{'{'{'b0,'bz,'b0xx0,'b0zz,'bz},'{'b1z0z,'bz,'b1zz,'b1zz,'b10z}},'{'{'bz,'b1xxzx,'b1xz,'bx0,'bzz1},'{'b1zz10,'bz,'bx,'b1,'b1x1z0}},'{'{'b0,'b0,'bzx11,'b0xz,'b010xx},'{'b1,'bzx1,'bz,'bz010,'b0z1}}},'{'{'{'b1,'b1,'bx0z,'b00x,'b1zx0},'{'b0x1z,'b001z,'b1xzx,'b0xz,'b00z}},'{'{'bx,'b01x11,'b11z1,'b1,'bxzzzz},'{'bz0,'bz,'b0zx,'b1xz,'bx}},'{'{'b0z,'b0,'bxzzx,'bz,'b0x},'{'bxz1x,'bzx,'b1z00,'b1,'b100x}}}};
  assign vwsbam = vwsbam;
endmodule: mf



// Seed after: 17955976471768091138,3128299129089410139
