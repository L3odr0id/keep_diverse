// Seed: 13809556470856728717,3128299129089410139

module ysbfobo
  ( output bit [1:4][2:4][4:3]  rio
  , output trireg logic [4:3][0:2][3:4] dcvacoxs [3:3][2:1][0:1]
  , output logic [3:1][4:3][4:3]  j
  , output wire logic [0:3][2:4][3:2][4:1] svrbcfg [1:2][2:3][4:2][1:3]
  , input shortreal tpr
  , input real ccjzwticew [1:0][4:1]
  );
  
  
  and qxad(jamineree, lkisy, g);
  
  not tfbl(xkb, dzooevekyp);
  
  not mrqegdzfk(j, eiez);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic j -> logic [3:1][4:3][4:3]  j
  
  
  // Single-driven assigns
  assign rio = '{'{'{'b0,'b0011},'{'b00,'b111},'{'b11,'b0}},'{'{'b0110,'b0100},'{'b11100,'b110},'{'b1000,'b1}},'{'{'b01,'b1},'{'b001,'b0001},'{'b1,'b00}},'{'{'b000,'b0010},'{'b10,'b000},'{'b0111,'b1000}}};
  
  // Multi-driven assigns
  assign eiez = lkisy;
endmodule: ysbfobo

module gkfezskbix
  ( output byte ottdunc [3:4]
  , output wor logic hvvoestrt [2:2]
  , output tri logic [2:2][1:3] h [2:3][0:0][3:2]
  , input triand logic [3:0] jnixbhnoxl [3:3][3:0][2:1][4:1]
  , input tri0 logic [2:3][3:4][2:3][3:4] tromr [3:0][1:1]
  );
  
  
  xor djkr(mhpbvyyl, zlrkqtigvd, xeamis);
  
  
  // Single-driven assigns
  assign ottdunc = ottdunc;
  
  // Multi-driven assigns
  assign h = h;
  assign xeamis = 'bxx1zx;
  assign zlrkqtigvd = 'bz101;
endmodule: gkfezskbix

module anbs
  ( output tri1 logic kko [0:4][3:3]
  , output bit baohsreh
  , output realtime grkct
  , output realtime vecbxfrfzs
  , input bit nqfrtrhfvo [1:4]
  , input triand logic atgyrg [2:4][2:2][3:3][3:2]
  , input logic [4:2][2:3][1:4]  t
  );
  
  
  not xisqyf(arfoyawf, baohsreh);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit baohsreh -> logic baohsreh
  
  
  // Single-driven assigns
  assign baohsreh = 'b101;
  assign grkct = baohsreh;
  
  // Multi-driven assigns
  assign kko = '{'{'b0x0zx},'{'b0z},'{'bxz},'{'b1z},'{'b0x}};
  assign arfoyawf = 'bz0x;
  assign atgyrg = '{'{'{'{'bz,'bzx0x}}},'{'{'{'b11x,'bx0x}}},'{'{'{'b101,'bx}}}};
endmodule: anbs



// Seed after: 9931058363952773939,3128299129089410139
