// Seed: 549568144774216018,3128299129089410139

module dhtgi
  (output tri1 logic [0:1][4:0][0:4] zqc [0:1], output shortreal kpjxhmfzhn, output shortreal wueuwijt);
  
  
  not ljuk(hju, kpjxhmfzhn);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal kpjxhmfzhn -> logic kpjxhmfzhn
  
  
  // Single-driven assigns
  assign kpjxhmfzhn = 'b0zzz0;
  
  // Multi-driven assigns
  assign zqc = '{'{'{'{'b111xx,'b11z,'b0x,'b11z10,'bxxx0x},'{'b1,'b0,'b1xzx1,'b1zzzx,'b01xxz},'{'b1101,'b0,'b100,'b1x00x,'b1xx1x},'{'b001,'b0,'bxz,'b1100,'b11z0x},'{'b00z,'bx11z,'bzz,'bz0,'b01000}},'{'{'b0zz,'b0,'b1z1x1,'bx,'b01},'{'b0z1,'bzxxx,'bz0z00,'b0,'b00xz},'{'b0010,'bx0xx,'bx1x0z,'b1z,'bz10zz},'{'b01zxx,'b11x1,'bx1,'b01,'bx00x},'{'bz,'bz,'b110,'b0x1,'bz}}},'{'{'{'b1zz,'bx0,'bzx,'b111x,'b0},'{'bzz,'bzx,'bx0z,'b1z0z,'b11},'{'b01x01,'bz0x01,'b0,'bxz1z,'b0100},'{'b0z,'bz1zxz,'b0011,'bx,'bzxzz1},'{'b0,'bx0,'bxx,'b011x0,'bzx0}},'{'{'bxx0z1,'bz,'bxxx,'b0,'b0xz0},'{'bxz1z0,'bzz1,'bz00z,'bz,'bz},'{'b11,'bz0000,'bz11,'b0x,'b1zx},'{'b0,'b1zxz,'bx1z1,'b1,'b1z1z0},'{'b0x,'b1z,'b1zz0,'b0,'b1xzz1}}}};
  assign hju = hju;
endmodule: dhtgi

module s
  ( output reg [2:0][0:2][2:2][3:2]  tdsp
  , output tri0 logic [3:0][4:2][4:3][1:3] knxuua [4:0]
  , output supply0 logic [4:2][3:3][0:1][0:2] tjyuq [4:1][1:3][4:1][0:0]
  , input wor logic [1:2][2:0][1:2][0:2] x [3:3][3:1][0:0][1:0]
  );
  
  
  not dbfzhoxvkv(tdsp, rgalgssik);
  // warning: implicit conversion of port connection expands from 1 to 18 bits
  //   logic tdsp -> reg [2:0][0:2][2:2][3:2]  tdsp
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign knxuua = knxuua;
  assign x = x;
  assign rgalgssik = rgalgssik;
  assign tjyuq = tjyuq;
endmodule: s

module dadcgeme
  ( output supply0 logic [4:0][0:1][1:0][3:1] mkgcbom [0:2]
  , output tri0 logic [1:2][4:3] grfoernyb [0:4][3:4][0:3]
  , output wand logic [3:4][0:1] gmkym [0:1]
  , output logic [1:4][4:1] hupqdyc [2:1]
  , input real gpnyi [0:1][1:0][4:2]
  , input uwire logic [3:2][3:2][3:0][2:1]  b
  );
  
  
  nand hpfszam(umhnduadao, n, xgfhqdyjdk);
  
  and clq(n, b, ouiu);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   uwire logic [3:2][3:2][3:0][2:1]  b -> logic b
  
  not ifhvegbn(beclonkmv, umhnduadao);
  
  not d(n, n);
  
  
  // Single-driven assigns
  assign hupqdyc = hupqdyc;
  
  // Multi-driven assigns
  assign mkgcbom = mkgcbom;
endmodule: dadcgeme



// Seed after: 9058340612855349718,3128299129089410139
