// Seed: 10476335463025953815,3128299129089410139

module yhdyae
  (output supply1 logic [3:2][3:0][2:2][2:1] kzmki [0:4][3:2][1:4], output uwire logic cabc, output logic [4:3][0:0] q [4:2]);
  
  
  not aavi(uxmzmksdmq, cabc);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kzmki = kzmki;
  assign uxmzmksdmq = 'b0x1z;
endmodule: yhdyae

module nwye
  ( output logic [1:4][4:0]  axgvat
  , output reg zhus
  , output supply0 logic [1:1]  ubtopvqr
  , output logic [1:1] woaznojn [1:1]
  , input shortint vhmnyqtsy
  , input bit [2:3]  ul
  , input wor logic [3:0][2:0][4:3][4:1] dejbxtytj [3:4][3:1][2:0]
  );
  
  logic [4:3][0:0] ao [4:2];
  supply1 logic [3:2][3:0][2:2][2:1] nuuoazkfpw [0:4][3:2][1:4];
  
  yhdyae mobagli(.kzmki(nuuoazkfpw), .cabc(axgvat), .q(ao));
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  //   uwire logic cabc -> logic [1:4][4:0]  axgvat
  
  not spgksujt(ubtopvqr, ul);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3]  ul -> logic ul
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ubtopvqr = vhmnyqtsy;
endmodule: nwye

module hjndgm
  ( output shortint dbrgtbv [3:2]
  , output tri logic [2:0][1:1] piiofi [2:0][0:2][3:2]
  , output wire logic [1:3][0:0][3:4] xd [2:4]
  , output tri logic [2:3]  qkhtkxydts
  , input wor logic ucgvohj
  , input wand logic [2:0] sl [1:4][3:3]
  , input logic [2:2][1:4][4:3]  unsxxugv
  , input reg [4:3][4:2][1:1]  rywsdeiprp
  );
  
  
  
  // Single-driven assigns
  assign dbrgtbv = dbrgtbv;
  
  // Multi-driven assigns
  assign qkhtkxydts = '{'bz0,'bzzxx};
endmodule: hjndgm

module lkjdgly
  (output logic hfwsyq [1:1][4:2][2:1][3:0], output bit rodb, output logic [0:1] dwb [3:1]);
  
  
  not shrmaq(rodb, rodb);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic rodb -> bit rodb
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit rodb -> logic rodb
  
  and jq(fvotwvmzf, rodb, aeueffuktf);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit rodb -> logic rodb
  
  not gbvnyvnugg(bhnr, lwlaoc);
  
  nand rdp(fvotwvmzf, fjhzqos, wtalkag);
  
  
  // Single-driven assigns
  assign hfwsyq = '{'{'{'{'b1x0zz,'b0xzx,'bzxxz0,'bz01x},'{'b1zzx,'bxz0,'b01011,'b10}},'{'{'b1xz,'bz10,'bxz0z,'bx},'{'bz1zx1,'b1,'b0zz,'bz}},'{'{'b1,'bx00z0,'bz0,'bz},'{'bzz,'bz,'bz,'b100}}}};
  
  // Multi-driven assigns
  assign wtalkag = 'b01111;
  assign lwlaoc = 'bx;
  assign fjhzqos = 'bzx11x;
  assign aeueffuktf = 'b0x0;
endmodule: lkjdgly



// Seed after: 8355443864916960300,3128299129089410139
