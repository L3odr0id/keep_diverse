// Seed: 7952459965154144426,3128299129089410139

module rcasvpw
  ( output uwire logic dsxvkecdmm
  , input reg [0:4][0:4] cigcb [2:3]
  , input wor logic tg [0:4][0:0][0:2]
  , input trireg logic kc [3:2]
  , input uwire logic stwhloq [4:0][3:0]
  );
  
  
  xor xphutwsae(yngvlbgj, k, dsxvkecdmm);
  
  and jxeajn(addrdvi, dsxvkecdmm, dsxvkecdmm);
  
  not iudjtyhogx(ju, hbdej);
  
  not u(lkqxvpek, lkqxvpek);
  
  
  // Single-driven assigns
  assign dsxvkecdmm = 'bx1x;
  
  // Multi-driven assigns
endmodule: rcasvpw

module piekw
  ( output tri0 logic [2:0][0:4][1:3] udz [1:3][1:4]
  , output trireg logic [0:4][1:2] ampvzzae [4:1][2:4][0:3][3:4]
  , output bit [2:2] nh [3:3]
  , output logic [4:1][0:1]  mkwvkbtat
  , input wire logic [0:0][0:1][3:0] tqwskncbg [1:2]
  );
  
  
  or gd(mkwvkbtat, vklum, vklum);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   logic mkwvkbtat -> logic [4:1][0:1]  mkwvkbtat
  
  or rugbzmfb(cbtclwu, ozffpvy, cbtclwu);
  
  
  // Single-driven assigns
  assign nh = nh;
  
  // Multi-driven assigns
  assign udz = udz;
endmodule: piekw



// Seed after: 15791412969388589653,3128299129089410139
