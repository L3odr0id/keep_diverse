// Seed: 3385037440923941020,3128299129089410139

module iudsxfwjem
  (output tri logic [2:0][2:0] ku [2:1][4:3], output reg [0:1][2:3] z [3:2], output wand logic yjdf [3:4][0:3]);
  
  
  or suujeuxccs(ff, ff, ff);
  
  xor gfjvozvny(enadcxhwj, ff, ntdjht);
  
  not la(wdud, btz);
  
  nand nmwvvelm(ff, ntdjht, jekwrkqfxs);
  
  
  // Single-driven assigns
  assign z = z;
  
  // Multi-driven assigns
  assign btz = 'bx1zx;
  assign ku = ku;
  assign ff = ff;
endmodule: iudsxfwjem

module kzzjrpgxin
  ( output tri0 logic [0:1]  thtyuvy
  , output tri1 logic [3:1][2:3] txxgjnh [2:3]
  , input reg [0:2][2:0][1:3]  mt
  , input logic [3:3][4:2][0:3] pjchanzsdm [2:3]
  );
  
  wand logic clzggfca [3:4][0:3];
  reg [0:1][2:3] cqgsssp [3:2];
  wand logic tehmevlvqz [3:4][0:3];
  reg [0:1][2:3] uuqtsekc [3:2];
  tri logic [2:0][2:0] lwt [2:1][4:3];
  
  iudsxfwjem kbrij(.ku(lwt), .z(uuqtsekc), .yjdf(tehmevlvqz));
  
  iudsxfwjem fwofuykaql(.ku(lwt), .z(cqgsssp), .yjdf(clzggfca));
  
  and lrcxqmbwml(thtyuvy, thtyuvy, thtyuvy);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic thtyuvy -> tri0 logic [0:1]  thtyuvy
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri0 logic [0:1]  thtyuvy -> logic thtyuvy
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri0 logic [0:1]  thtyuvy -> logic thtyuvy
  
  not xadmhsev(zqqorchae, thtyuvy);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri0 logic [0:1]  thtyuvy -> logic thtyuvy
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign clzggfca = tehmevlvqz;
  assign tehmevlvqz = '{'{'b0x,'b0x00x,'bz1x0,'bx0xz0},'{'b10,'b0,'b10zx,'bzzz}};
  assign thtyuvy = thtyuvy;
endmodule: kzzjrpgxin



// Seed after: 8966281038822525192,3128299129089410139
