// Seed: 5879450806462840495,3128299129089410139

module zuokjh
  ( output reg [3:3][4:2][0:3]  qvr
  , output bit [1:1]  vsdcwlmsvh
  , output reg [1:0] vaq [4:3][2:4]
  , output tri logic [1:3][2:0][0:1] qw [4:2][2:1][2:3]
  , input byte gm
  );
  
  
  and impkz(ts, qvr, qvr);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [3:3][4:2][0:3]  qvr -> logic qvr
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [3:3][4:2][0:3]  qvr -> logic qvr
  
  xor uqqzsierx(bgsywz, gm, quxtxlt);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte gm -> logic gm
  
  nand j(dyrcnwi, wpuu, qogxmsien);
  
  
  // Single-driven assigns
  assign qvr = vsdcwlmsvh;
  
  // Multi-driven assigns
  assign bgsywz = vsdcwlmsvh;
endmodule: zuokjh

module chdpghefof
  ( output supply0 logic [2:3][0:0][0:1][0:2] dmpxkgemy [0:2][2:1][4:3]
  , input tri logic [2:0][3:2][0:1] cvlqnwhv [1:3][3:2]
  , input reg [2:3][2:3][0:2]  pmzkkm
  );
  
  
  or rbvlv(ptmwztsb, ptmwztsb, ptmwztsb);
  
  not cwd(jubmyyb, ptmwztsb);
  
  and up(ppgcofrkb, ptmwztsb, n);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign n = 'bxxx;
  assign dmpxkgemy = dmpxkgemy;
  assign ptmwztsb = 'b0zz;
endmodule: chdpghefof



// Seed after: 12475482197253238135,3128299129089410139
