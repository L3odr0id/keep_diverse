// Seed: 16610296227259165878,3128299129089410139

module iwcnxgowym
  (output reg [2:2][1:4]  wf, output reg [3:4][1:0][3:2]  sgigakm);
  
  
  xor fjcp(kbonxtex, qyijvy, hjebzwiiwk);
  
  or evt(wf, msy, kayd);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic wf -> reg [2:2][1:4]  wf
  
  not apvqgwykud(uy, wf);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   reg [2:2][1:4]  wf -> logic wf
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kayd = 'b00;
  assign kbonxtex = wf;
endmodule: iwcnxgowym

module emfqvezkoa
  ( output tri0 logic [1:2][3:3] ldhyk [3:2][3:3]
  , output time j [1:4][2:1][2:4]
  , output logic pjl
  , output time ukya
  , input supply1 logic [2:4][4:3][3:4][3:2] zimivj [2:3][0:3][0:4][1:1]
  , input bit [0:4][0:3]  z
  );
  
  
  xor x(okmprgfbt, pjl, z);
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:4][0:3]  z -> logic z
  
  
  // Single-driven assigns
  assign j = '{'{'{'b1zx,'bzx1z,'bz00z},'{'bz11x1,'b111x,'b0xz}},'{'{'b10,'b1,'b1},'{'bxz0,'bz101,'bxxz}},'{'{'bzz011,'b101x,'b1},'{'bzz,'b000,'b010}},'{'{'bx0zx1,'b1xxxz,'bxz},'{'b0x1x,'bx0x,'b0110}}};
  
  // Multi-driven assigns
endmodule: emfqvezkoa



// Seed after: 16247055769448328577,3128299129089410139
