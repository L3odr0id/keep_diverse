// Seed: 1276793512140722276,3128299129089410139

module qxdqmrx
  ( output triand logic [3:1][3:1][4:2]  demltpbhiz
  , output bit [2:4][1:3][2:4]  wm
  , output supply0 logic [2:3] dyu [1:1][4:1]
  , output wire logic [2:2][3:2][2:3] kuerqyau [3:3][4:1]
  , input reg [1:4][4:1][3:2]  nllwipcvgy
  , input real demymn
  , input supply0 logic gzalucvbu [4:4][3:4][0:3][2:0]
  , input tri0 logic [3:0][3:4] hcuftfkg [1:4][1:4]
  );
  
  
  and hazh(grrmbja, wm, demymn);
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][1:3][2:4]  wm -> logic wm
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real demymn -> logic demymn
  
  not s(erjcfbb, xjkpx);
  
  not ejz(demltpbhiz, xjkpx);
  // warning: implicit conversion of port connection expands from 1 to 27 bits
  //   logic demltpbhiz -> triand logic [3:1][3:1][4:2]  demltpbhiz
  
  and rrk(twjlkvev, demltpbhiz, mlphsl);
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  //   triand logic [3:1][3:1][4:2]  demltpbhiz -> logic demltpbhiz
  
  
  // Single-driven assigns
  assign wm = demltpbhiz;
  
  // Multi-driven assigns
endmodule: qxdqmrx

module ydzugbnr
  ( output reg v [0:1][2:3]
  , output tri1 logic [0:2][4:2][4:4] gbml [0:3][2:1]
  , output byte pjjrlr [4:4]
  , input wire logic [0:2] si [0:0][4:1][2:0][1:0]
  , input real ijkow
  , input wire logic kzylgfudt [3:0][1:4][1:3][0:1]
  );
  
  
  not cg(u, gqg);
  
  
  // Single-driven assigns
  assign v = v;
  
  // Multi-driven assigns
  assign gqg = u;
  assign gbml = gbml;
endmodule: ydzugbnr

module imbtvb
  (input supply0 logic [3:3][1:3]  cpq, input logic [2:4][3:2] x [1:3][3:0]);
  
  wire logic [2:2][3:2][2:3] mellxvtk [3:3][4:1];
  supply0 logic [2:3] jg [1:1][4:1];
  tri0 logic [3:0][3:4] ydnbcqbgk [1:4][1:4];
  supply0 logic pp [4:4][3:4][0:3][2:0];
  
  qxdqmrx t(.demltpbhiz(yszle), .wm(cpq), .dyu(jg), .kuerqyau(mellxvtk), .nllwipcvgy(cpq), .demymn(cpq), .gzalucvbu(pp), .hcuftfkg(ydnbcqbgk));
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  //   triand logic [3:1][3:1][4:2]  demltpbhiz -> wire logic yszle
  //
  // warning: implicit conversion of port connection truncates from 27 to 3 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][1:3][2:4]  wm -> supply0 logic [3:3][1:3]  cpq
  //
  // warning: implicit conversion of port connection expands from 3 to 32 bits
  //   supply0 logic [3:3][1:3]  cpq -> reg [1:4][4:1][3:2]  nllwipcvgy
  //
  // warning: implicit conversion of port connection expands from 3 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   supply0 logic [3:3][1:3]  cpq -> real demymn
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign cpq = '{'{'bx110,'bxx,'bxxxz}};
  assign ydnbcqbgk = '{'{'{'{'bx1,'bzx},'{'b1,'bz00},'{'b0zx1,'b0xz},'{'bzzzxx,'b10x}},'{'{'bz01z1,'b1},'{'bxx0xx,'bxz},'{'b0xxx,'b0x0},'{'bz1,'b00}},'{'{'bzxxz1,'bz1},'{'b01,'bzx},'{'bxzxz0,'b010},'{'bz,'bxz00}},'{'{'bzxxxz,'b0xzz1},'{'b1z1z,'bz0xz},'{'b0x1x1,'bx0z1},'{'b101x,'bxz1x}}},'{'{'{'b1,'b1000},'{'b1z101,'b1zx},'{'bz,'bx},'{'b1xx,'b0x0z}},'{'{'b0,'b0x0zx},'{'b1,'b10x},'{'bx0,'bx1z},'{'b111x,'b1x100}},'{'{'bx,'bz},'{'b1zz1z,'bx0x1},'{'b0z0,'bz},'{'bz,'b1x1}},'{'{'b0xxx,'b00zxz},'{'b1xz,'b01},'{'b011,'bx},'{'bx0x01,'bxz01z}}},'{'{'{'bz111x,'bzxz},'{'bz0zx0,'bzx},'{'b00,'b10zz1},'{'bxx,'bxzz1}},'{'{'bx01x,'bzxzz},'{'bzzx,'b1xxz0},'{'bz,'b1zz},'{'bx010x,'b0}},'{'{'bx,'b0zx},'{'bz,'bx1z1},'{'bz00,'bxxx1},'{'bzx10,'b1x0}},'{'{'b100zz,'bx},'{'bx1xx,'b0z00},'{'bz1,'b11z},'{'bz0zxx,'b1}}},'{'{'{'bz,'b10zz0},'{'b1zz0,'bz},'{'b01x11,'b00x},'{'bz,'bxxz}},'{'{'bx0x1,'bxx0},'{'b0zz0,'bz},'{'b00xxx,'bx1zx0},'{'b00zxx,'bxzzx}},'{'{'b1,'b0x10},'{'bz0z11,'b1},'{'b1zzxz,'bx0},'{'bz,'b1z000}},'{'{'bzx,'bz1},'{'bz1x0z,'bx1zzx},'{'b101,'bx0},'{'b10,'bx}}}};
  assign pp = '{'{'{'{'b10z1,'bz,'b0},'{'bzzxx,'bz,'b101z},'{'b11x,'bzzx,'bzxz},'{'bz,'b00z00,'b0}},'{'{'b100zz,'bzz0,'b1xx1z},'{'bxz,'bz110,'b100},'{'bx1,'b00,'b1z1z},'{'bz,'bx,'bz}}}};
endmodule: imbtvb



// Seed after: 11378901856138186289,3128299129089410139
