// Seed: 14390351302887849332,3128299129089410139

module myhooo
  ( output bit [0:3] l [0:3][0:1][2:0]
  , input wand logic [0:2][2:3] apvi [1:0]
  , input reg [4:2][2:1][0:1] ymezhbzy [4:4]
  , input trireg logic [2:3][1:1] fwsjrkogju [2:2][4:1][4:3][2:2]
  , input tri logic ko [1:0][3:3][2:1]
  );
  
  
  not xkbvaq(vlylkx, kxieugldwl);
  
  nand ykwmusbacd(ist, iwzvbtra, ist);
  
  not vtpbgdunvd(les, otonkx);
  
  
  // Single-driven assigns
  assign l = '{'{'{'{'b1110,'b1000,'b11,'b00},'{'b1,'b00,'b0110,'b10},'{'b01,'b100,'b00,'b1}},'{'{'b1000,'b01,'b01,'b101},'{'b101,'b10100,'b0111,'b1},'{'b01111,'b00,'b11,'b1111}}},'{'{'{'b10,'b0,'b0,'b0111},'{'b01,'b01,'b10100,'b10100},'{'b101,'b0001,'b11,'b11}},'{'{'b1,'b1101,'b01,'b0111},'{'b00000,'b11,'b10,'b1},'{'b10,'b100,'b100,'b11100}}},'{'{'{'b111,'b0100,'b1,'b00},'{'b1110,'b11,'b0,'b11},'{'b00100,'b1,'b1101,'b0001}},'{'{'b10110,'b00,'b11000,'b1100},'{'b1,'b11,'b000,'b010},'{'b100,'b111,'b001,'b11}}},'{'{'{'b010,'b1101,'b000,'b0011},'{'b110,'b11100,'b10,'b10},'{'b01,'b010,'b1100,'b1111}},'{'{'b0000,'b01,'b1,'b00100},'{'b011,'b00,'b001,'b1},'{'b1,'b110,'b0110,'b10}}}};
  
  // Multi-driven assigns
  assign apvi = apvi;
  assign kxieugldwl = kxieugldwl;
endmodule: myhooo



// Seed after: 2189224357496412630,3128299129089410139
