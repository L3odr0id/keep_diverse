// Seed: 10452617400833083778,3128299129089410139

module xxgnjsjsp
  ( output int aczu
  , output triand logic [1:0][1:2][2:0] oiiqzdvo [1:4][1:3][4:3]
  , input logic uwqjv
  , input trireg logic hvamh [1:0][3:4]
  );
  
  
  
  // Single-driven assigns
  assign aczu = aczu;
  
  // Multi-driven assigns
  assign oiiqzdvo = oiiqzdvo;
  assign hvamh = '{'{'b1z01,'b00},'{'bx1xz,'b0zx1}};
endmodule: xxgnjsjsp



// Seed after: 10476335463025953815,3128299129089410139
