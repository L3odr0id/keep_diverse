// Seed: 5762705560976339521,3128299129089410139

module nwxdqo
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: nwxdqo

module abxcpm
  ( output tri logic [2:1][3:0] xjtsbu [1:4][0:4]
  , output tri logic [3:1][3:3][4:1][3:3] g [1:2][2:2][3:1][0:1]
  , input supply1 logic [2:0] b [3:3][4:3][1:3][4:3]
  , input int jmxtq [0:3][2:0]
  , input wire logic [0:0]  zwx
  );
  
  
  not yxgql(zwx, zwx);
  
  not ilcqppgxh(opqji, zwx);
  
  nwxdqo bnmu();
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: abxcpm

module yslksythrb
  ( output tri0 logic [2:1][4:0][0:1]  qnnzhmb
  , input real znwr
  , input realtime wavnisainn [3:4]
  , input bit [4:3][2:0][0:4]  ky
  , input bit qb [2:4]
  );
  
  tri logic [3:1][3:3][4:1][3:3] tor [1:2][2:2][3:1][0:1];
  tri logic [2:1][3:0] lzekdf [1:4][0:4];
  tri logic [3:1][3:3][4:1][3:3] wvnukhlie [1:2][2:2][3:1][0:1];
  tri logic [3:1][3:3][4:1][3:3] ih [1:2][2:2][3:1][0:1];
  tri logic [2:1][3:0] kzicevg [1:4][0:4];
  int m [0:3][2:0];
  supply1 logic [2:0] d [3:3][4:3][1:3][4:3];
  int pihntjvm [0:3][2:0];
  int burde [0:3][2:0];
  supply1 logic [2:0] y [3:3][4:3][1:3][4:3];
  
  abxcpm zeymss(.xjtsbu(kzicevg), .g(ih), .b(y), .jmxtq(burde), .zwx(qnnzhmb));
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   tri0 logic [2:1][4:0][0:1]  qnnzhmb -> wire logic [0:0]  zwx
  
  not ydvdw(qnnzhmb, kuspc);
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  //   logic qnnzhmb -> tri0 logic [2:1][4:0][0:1]  qnnzhmb
  
  abxcpm rfuvazud(.xjtsbu(kzicevg), .g(wvnukhlie), .b(y), .jmxtq(pihntjvm), .zwx(kuspc));
  
  abxcpm prw(.xjtsbu(lzekdf), .g(tor), .b(d), .jmxtq(m), .zwx(qnnzhmb));
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   tri0 logic [2:1][4:0][0:1]  qnnzhmb -> wire logic [0:0]  zwx
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: yslksythrb

module lshooa
  (output shortreal aszsul, input tri1 logic yyralitbc [0:3][3:1][3:0][2:3]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign yyralitbc = '{'{'{'{'b0x11,'b0100},'{'b0xz10,'b10xxx},'{'b0z1z1,'b1},'{'bx,'b0z10}},'{'{'bxz01,'bx},'{'bzx1,'bx},'{'b0,'bz},'{'b10,'bz}},'{'{'b1011,'b010z},'{'b1zzzz,'b1},'{'bx,'b1z0xz},'{'b010x,'b1z0zx}}},'{'{'{'bxx0x,'bx11},'{'bz,'b01},'{'bz01x,'b000},'{'bxxxx0,'b0x}},'{'{'b1,'bx},'{'bx001,'b01z},'{'bx1z,'b0x0},'{'bzx0,'bz}},'{'{'b1,'b10x},'{'bzz1zx,'bxz},'{'b1,'bx},'{'b1,'bz1x0}}},'{'{'{'bx0,'b111x},'{'bzz,'b1},'{'bzxxxx,'b0},'{'bx1011,'b110}},'{'{'bz0z,'bz0x01},'{'bx,'bxz10x},'{'bxzx01,'b01},'{'b1z,'bx0zx}},'{'{'bxzz,'b0111z},'{'bx0z1,'b0z},'{'b1,'b00},'{'b0z,'bxx}}},'{'{'{'b01z1,'b1x1},'{'bz11x1,'b1},'{'bz,'bx1zx},'{'b1,'b0x10}},'{'{'b000,'b0z},'{'bx01,'bx},'{'bx1,'bzzx},'{'b1x,'b11}},'{'{'bzz1,'b01x},'{'bx11z,'b1},'{'bxz0x,'bx},'{'b111,'b011xz}}}};
endmodule: lshooa



// Seed after: 5879450806462840495,3128299129089410139
