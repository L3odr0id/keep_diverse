// Seed: 11767764356932420300,3128299129089410139

module zioylimvij
  ( output longint s [3:0][2:4][3:0]
  , output tri1 logic [3:2][2:1][0:3][2:3] ind [4:2][0:2][4:4]
  , input tri logic [4:2] carngr [2:2]
  );
  
  
  nand zce(zchdmou, bhfhfn, bhfhfn);
  
  nand ensmnj(bhfhfn, bhfhfn, yi);
  
  not zpt(bhfhfn, bhfhfn);
  
  
  // Single-driven assigns
  assign s = s;
  
  // Multi-driven assigns
  assign ind = ind;
endmodule: zioylimvij



// Seed after: 2769780858164702270,3128299129089410139
