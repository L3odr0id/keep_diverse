// Seed: 328071024425920796,3128299129089410139

module baxg
  ( output uwire logic zy [2:3]
  , input logic [0:1]  ghdjrqo
  , input supply1 logic [3:0] nvf [3:1][2:3][3:2][1:4]
  , input tri logic [3:1][2:4][3:0][1:3] vnirwrxeq [4:4][1:0][4:4]
  , input realtime w [1:4][0:3]
  );
  
  
  not iwoxb(oeqzbhlxsn, oeqzbhlxsn);
  
  nand vxo(sspfdmhz, ir, oeqzbhlxsn);
  
  not mzddm(oeqzbhlxsn, sdxizgzti);
  
  nand rwquzzjsi(oeqzbhlxsn, ir, xa);
  
  
  // Single-driven assigns
  assign zy = '{'bxxx0x,'b1z};
  
  // Multi-driven assigns
  assign oeqzbhlxsn = ir;
  assign vnirwrxeq = vnirwrxeq;
endmodule: baxg

module qmr
  (output bit [4:4][0:0] ojtnbiqhjw [3:4][1:4], input tri0 logic [3:3][0:3][1:0] chayjfmeb [3:0]);
  
  uwire logic uiczhagc [2:3];
  realtime moyhmpbbv [1:4][0:3];
  tri logic [3:1][2:4][3:0][1:3] f [4:4][1:0][4:4];
  supply1 logic [3:0] szfkcbmhnw [3:1][2:3][3:2][1:4];
  
  baxg skr(.zy(uiczhagc), .ghdjrqo(fnrc), .nvf(szfkcbmhnw), .vnirwrxeq(f), .w(moyhmpbbv));
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   wire logic fnrc -> logic [0:1]  ghdjrqo
  
  or brdutydndl(fnrc, fnrc, fnrc);
  
  
  // Single-driven assigns
  assign ojtnbiqhjw = ojtnbiqhjw;
  assign moyhmpbbv = '{'{'bx0z00,'bx1x,'b010z,'bx11z},'{'b011z,'b0,'b101,'b0xz},'{'b1zz10,'bx11x0,'b1,'bxz0},'{'bz,'b00x0x,'bx,'b01}};
  
  // Multi-driven assigns
  assign fnrc = 'b101;
endmodule: qmr

module zye
  (output wand logic [2:0]  lvf, output tri1 logic [1:1]  pcgef, input shortint tcnt);
  
  
  not erzty(l, tcnt);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint tcnt -> logic tcnt
  
  and fqlbnmcgvz(aqj, duzrqznhy, lvf);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wand logic [2:0]  lvf -> logic lvf
  
  or ekmwywm(afwbk, bkoqyob, fszrtqkrgl);
  
  not dglc(qlpkzosfuz, jcclzmva);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign lvf = '{'bxz01z,'b1,'bx1z0};
  assign duzrqznhy = lvf;
endmodule: zye



// Seed after: 3969165351885200449,3128299129089410139
