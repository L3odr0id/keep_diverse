// Seed: 9947113201368221206,3128299129089410139

module vv
  (output triand logic [0:3][0:1][1:4][3:3] uxtvttw [0:0][4:2][2:4][1:0], output tri logic [1:0][3:3][3:1][4:0]  mcgiwhgfet, input reg cyduengbv);
  
  
  not ddxzuojim(mcgiwhgfet, mcgiwhgfet);
  // warning: implicit conversion of port connection expands from 1 to 30 bits
  //   logic mcgiwhgfet -> tri logic [1:0][3:3][3:1][4:0]  mcgiwhgfet
  //
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   tri logic [1:0][3:3][3:1][4:0]  mcgiwhgfet -> logic mcgiwhgfet
  
  not vjq(mcgiwhgfet, cyduengbv);
  // warning: implicit conversion of port connection expands from 1 to 30 bits
  //   logic mcgiwhgfet -> tri logic [1:0][3:3][3:1][4:0]  mcgiwhgfet
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign uxtvttw = uxtvttw;
  assign mcgiwhgfet = '{'{'{'{'b0z,'b0,'bz0x0,'b11,'b1z1xz},'{'bz10x0,'b1zx1z,'bzz1x,'bzxx,'bx1x1},'{'bz,'bz0,'b01011,'b10x,'b10z0}}},'{'{'{'b00z,'bxzzx,'b1011x,'b11xzz,'b1xz11},'{'b01,'bx1zz0,'bzx0z,'b1z,'bz01},'{'b10x,'bxx0z,'b111,'b0z0z1,'bxz0xx}}}};
endmodule: vv

module hpphm
  (input byte rhdmtlfblp, input reg vzjv, input reg [1:3][0:3][0:2]  alrutgvh, input trireg logic hh [3:1]);
  
  triand logic [0:3][0:1][1:4][3:3] wbppuht [0:0][4:2][2:4][1:0];
  
  vv vujmnt(.uxtvttw(wbppuht), .mcgiwhgfet(azttg), .cyduengbv(rhdmtlfblp));
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   tri logic [1:0][3:3][3:1][4:0]  mcgiwhgfet -> wire logic azttg
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte rhdmtlfblp -> reg cyduengbv
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign wbppuht = wbppuht;
  assign hh = '{'b10,'b01,'bz11};
endmodule: hpphm

module rhiovc
  ( output reg [1:1][4:2][0:1]  kvvsdt
  , output bit [3:1] hjqp [1:2]
  , output reg [0:1] ws [0:1][1:1]
  , input supply0 logic [4:2] dyrz [0:2][4:3][3:0][2:3]
  , input tri0 logic [2:1][2:2][2:4][3:2] ljpcsl [2:4][3:1][0:2]
  , input logic [0:0][3:3]  afjsxmb
  );
  
  
  and nwgt(kvvsdt, afjsxmb, rbfyowxie);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   logic kvvsdt -> reg [1:1][4:2][0:1]  kvvsdt
  
  or gse(dij, rbfyowxie, dij);
  
  
  // Single-driven assigns
  assign ws = ws;
  assign hjqp = '{'{'b1,'b0,'b0110},'{'b1111,'b11100,'b0}};
  
  // Multi-driven assigns
endmodule: rhiovc



// Seed after: 1735739043436887574,3128299129089410139
