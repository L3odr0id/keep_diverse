// Seed: 1148233422042294380,3128299129089410139

module daoiggc
  ( output real zlcbqjpw [2:4][1:1]
  , output shortreal uvrxgmq
  , output bit [4:2]  xktwai
  , output triand logic [1:4][0:3] jkpkl [2:4][0:1]
  , input int newegrwuem [4:3][3:2]
  , input tri logic [1:3] bt [2:4]
  , input reg [4:3][0:2]  crxuuxoh
  , input uwire logic [2:2][2:1] vsmses [4:4][0:3]
  );
  
  
  not asbcyf(uvrxgmq, uvrxgmq);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic uvrxgmq -> shortreal uvrxgmq
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal uvrxgmq -> logic uvrxgmq
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jkpkl = jkpkl;
  assign bt = bt;
endmodule: daoiggc



// Seed after: 549568144774216018,3128299129089410139
