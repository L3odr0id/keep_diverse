// Seed: 16301470472216710936,3128299129089410139

module okr
  ( input triand logic cvfrzlew
  , input logic [2:3][3:2] rz [0:2]
  , input supply1 logic [1:2][1:2] ziaaqr [0:3][0:2][3:0]
  , input trireg logic [3:2][0:2]  oyqkv
  );
  
  
  or cpqacyqyp(oyqkv, oyqkv, oyqkv);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   logic oyqkv -> trireg logic [3:2][0:2]  oyqkv
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   trireg logic [3:2][0:2]  oyqkv -> logic oyqkv
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   trireg logic [3:2][0:2]  oyqkv -> logic oyqkv
  
  not qqngny(oyqkv, cvfrzlew);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   logic oyqkv -> trireg logic [3:2][0:2]  oyqkv
  
  nand uuoam(oyqkv, cvfrzlew, k);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   logic oyqkv -> trireg logic [3:2][0:2]  oyqkv
  
  not s(k, oyqkv);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   trireg logic [3:2][0:2]  oyqkv -> logic oyqkv
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign oyqkv = cvfrzlew;
  assign cvfrzlew = 'bzx10x;
endmodule: okr



// Seed after: 15923648016595859751,3128299129089410139
