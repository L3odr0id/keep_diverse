// Seed: 16536538239648392389,3128299129089410139

module er
  ( output logic ublsinf [0:2]
  , output uwire logic [4:4][0:4] ov [0:2][1:3][2:0][4:1]
  , output supply1 logic [4:4] ovyuktg [1:1]
  , output logic [0:1][2:2]  tjdziw
  , input wand logic [3:1][0:4] nxyzsf [1:2][3:0]
  , input shortreal yzeyaejymx
  , input logic qihjsjhw
  , input logic [3:4]  g
  );
  
  
  not biilrdc(tjdziw, g);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic tjdziw -> logic [0:1][2:2]  tjdziw
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [3:4]  g -> logic g
  
  xor ozxkvgow(vfpfymjl, ksjtzh, hee);
  
  xor iuvvavza(fxf, vfpfymjl, tjdziw);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [0:1][2:2]  tjdziw -> logic tjdziw
  
  nand fqc(ksjtzh, ksjtzh, qihjsjhw);
  
  
  // Single-driven assigns
  assign ublsinf = ublsinf;
  assign ov = ov;
  
  // Multi-driven assigns
  assign hee = tjdziw;
  assign ovyuktg = ovyuktg;
endmodule: er



// Seed after: 10931487316550548278,3128299129089410139
