// Seed: 4427233426964322947,3128299129089410139

module haidfe
  (output bit [3:3] dqoy [1:0][3:1]);
  
  
  not wxqgawmor(fwbpxhwe, o);
  
  or egenddntgd(yklxxsmvy, o, vqgksw);
  
  
  // Single-driven assigns
  assign dqoy = '{'{'{'b00001},'{'b0},'{'b100}},'{'{'b0010},'{'b1110},'{'b001}}};
  
  // Multi-driven assigns
endmodule: haidfe



// Seed after: 3385037440923941020,3128299129089410139
