// Seed: 14973839198957523227,3128299129089410139

module ded
  (output logic [3:2][1:3][0:3]  kiywmkuqs, output tri logic [2:1][0:2]  pfoo, output supply0 logic twgpjtikfk [4:0]);
  
  
  not bza(kiywmkuqs, kiywmkuqs);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic kiywmkuqs -> logic [3:2][1:3][0:3]  kiywmkuqs
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   logic [3:2][1:3][0:3]  kiywmkuqs -> logic kiywmkuqs
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ded

module vqrbmcnmq
  ( output wand logic [0:0][2:1] t [2:4]
  , output wire logic ppm [3:1][0:0][2:2]
  , output tri logic [3:1][1:1][4:1][2:3] lee [1:1]
  , output logic [0:3][1:4]  fdpfitugc
  );
  
  
  not wzn(dupc, ynrjqcb);
  
  
  // Single-driven assigns
  assign fdpfitugc = '{'{'bz0,'b0z1,'bz0xx,'bz0z1x},'{'b1x0,'bx01,'bxx,'b1z11z},'{'b10,'b0z0,'b1,'bx1zx},'{'bx,'bx0011,'b00,'b0z}};
  
  // Multi-driven assigns
  assign dupc = 'b0x1;
  assign lee = lee;
  assign ppm = '{'{'{'b0x0z}},'{'{'b1x}},'{'{'bxz0}}};
  assign t = '{'{'{'bxx111,'bx}},'{'{'b0011,'b01001}},'{'{'b01z10,'bz0z0}}};
endmodule: vqrbmcnmq

module uorufjcqa
  (output reg [1:2][0:3][2:3][4:3]  sfy, input supply1 logic fjtr [2:1][3:3][3:3][3:1]);
  
  
  
  // Single-driven assigns
  assign sfy = sfy;
  
  // Multi-driven assigns
  assign fjtr = fjtr;
endmodule: uorufjcqa

module axzfvplqc
  ( output realtime xz [2:3][4:2][4:4]
  , output logic [0:3][4:1][0:4][0:2]  zyikrdwls
  , output trireg logic [0:4] ciagq [2:1]
  , input uwire logic [2:2][1:1] vqfwm [3:4][0:0]
  , input reg htakqcpmjo [4:1]
  , input bit [0:1][1:1]  vcdxyjdy
  , input bit [3:2][4:1][4:2][1:3]  rnlwqcba
  );
  
  
  not mmcnccpxka(zyikrdwls, vcdxyjdy);
  // warning: implicit conversion of port connection expands from 1 to 240 bits
  //   logic zyikrdwls -> logic [0:3][4:1][0:4][0:2]  zyikrdwls
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:1][1:1]  vcdxyjdy -> logic vcdxyjdy
  
  
  // Single-driven assigns
  assign xz = xz;
  
  // Multi-driven assigns
  assign ciagq = ciagq;
endmodule: axzfvplqc



// Seed after: 7952459965154144426,3128299129089410139
