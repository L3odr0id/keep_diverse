// Seed: 2519640146387862472,3128299129089410139

module tejrmeyozf
  ( output integer qhnrulfyhu
  , output wor logic [0:1][1:2][1:4]  pbbplpwym
  , output wor logic [3:2][0:3][1:4]  vfvnsb
  , output shortreal gvtn [2:0][0:1]
  , input tri logic [1:2] axjjou [0:0][0:3][2:2]
  );
  
  
  
  // Single-driven assigns
  assign qhnrulfyhu = pbbplpwym;
  
  // Multi-driven assigns
  assign pbbplpwym = '{'{'{'b1zzx,'b1z001,'bxx,'b0zz},'{'bz0,'b101zz,'bxx,'bx0x0}},'{'{'bx,'bx,'b00x0z,'b1001},'{'b0x0,'b0xx1,'b0,'bx}}};
  assign axjjou = axjjou;
  assign vfvnsb = '{'{'{'b101,'bx0zx,'bzz,'b11100},'{'bz,'bz0,'bzz00x,'bz00z},'{'bxz10,'b1xx,'b1z,'b0xz1},'{'bx0101,'b0,'b10x0,'b1x0}},'{'{'bz,'bz,'bx,'bx},'{'bx0,'bxxz0,'bxx0,'b1z1},'{'bz11x,'bz,'b0z000,'b10},'{'b1x,'bxxx,'b111,'b0}}};
endmodule: tejrmeyozf



// Seed after: 2461222892141417034,3128299129089410139
